magic
tech sky130A
timestamp 1722865417
<< error_p >>
rect 150 2100 350 2550
<< dnwell >>
rect 150 1995 455 4055
<< nwell >>
rect 150 3950 500 4850
rect 350 2100 500 3950
rect 150 1200 500 2100
<< pwell >>
rect 200 3850 300 3900
rect 250 2200 300 3850
rect 200 2150 300 2200
<< psubdiff >>
rect 200 4935 600 4950
rect 200 4915 215 4935
rect 235 4915 265 4935
rect 285 4915 315 4935
rect 335 4915 365 4935
rect 385 4915 415 4935
rect 435 4915 465 4935
rect 485 4915 515 4935
rect 535 4915 565 4935
rect 585 4915 600 4935
rect 200 4900 600 4915
rect 550 4885 600 4900
rect 550 4865 565 4885
rect 585 4865 600 4885
rect 550 4835 600 4865
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 200 3885 300 3900
rect 200 3865 215 3885
rect 235 3865 265 3885
rect 285 3865 300 3885
rect 200 3850 300 3865
rect 250 3835 300 3850
rect 250 3815 265 3835
rect 285 3815 300 3835
rect 250 3785 300 3815
rect 250 3765 265 3785
rect 285 3765 300 3785
rect 250 3735 300 3765
rect 250 3715 265 3735
rect 285 3715 300 3735
rect 250 3685 300 3715
rect 250 3665 265 3685
rect 285 3665 300 3685
rect 250 3635 300 3665
rect 250 3615 265 3635
rect 285 3615 300 3635
rect 250 3585 300 3615
rect 250 3565 265 3585
rect 285 3565 300 3585
rect 250 3535 300 3565
rect 250 3515 265 3535
rect 285 3515 300 3535
rect 250 3485 300 3515
rect 250 3465 265 3485
rect 285 3465 300 3485
rect 250 3435 300 3465
rect 250 3415 265 3435
rect 285 3415 300 3435
rect 250 3385 300 3415
rect 250 3365 265 3385
rect 285 3365 300 3385
rect 250 3335 300 3365
rect 250 3315 265 3335
rect 285 3315 300 3335
rect 250 3285 300 3315
rect 250 3265 265 3285
rect 285 3265 300 3285
rect 250 3235 300 3265
rect 250 3215 265 3235
rect 285 3215 300 3235
rect 250 3185 300 3215
rect 250 3165 265 3185
rect 285 3165 300 3185
rect 250 3135 300 3165
rect 250 3115 265 3135
rect 285 3115 300 3135
rect 250 3085 300 3115
rect 250 3065 265 3085
rect 285 3065 300 3085
rect 250 3035 300 3065
rect 250 3015 265 3035
rect 285 3015 300 3035
rect 250 2985 300 3015
rect 250 2965 265 2985
rect 285 2965 300 2985
rect 250 2935 300 2965
rect 250 2915 265 2935
rect 285 2915 300 2935
rect 250 2885 300 2915
rect 250 2865 265 2885
rect 285 2865 300 2885
rect 250 2835 300 2865
rect 250 2815 265 2835
rect 285 2815 300 2835
rect 250 2785 300 2815
rect 250 2765 265 2785
rect 285 2765 300 2785
rect 250 2735 300 2765
rect 250 2715 265 2735
rect 285 2715 300 2735
rect 250 2685 300 2715
rect 250 2665 265 2685
rect 285 2665 300 2685
rect 250 2635 300 2665
rect 250 2615 265 2635
rect 285 2615 300 2635
rect 250 2585 300 2615
rect 250 2565 265 2585
rect 285 2565 300 2585
rect 250 2535 300 2565
rect 250 2515 265 2535
rect 285 2515 300 2535
rect 250 2485 300 2515
rect 250 2465 265 2485
rect 285 2465 300 2485
rect 250 2435 300 2465
rect 250 2415 265 2435
rect 285 2415 300 2435
rect 250 2385 300 2415
rect 250 2365 265 2385
rect 285 2365 300 2385
rect 250 2335 300 2365
rect 250 2315 265 2335
rect 285 2315 300 2335
rect 250 2285 300 2315
rect 250 2265 265 2285
rect 285 2265 300 2285
rect 250 2235 300 2265
rect 250 2215 265 2235
rect 285 2215 300 2235
rect 250 2200 300 2215
rect 200 2185 300 2200
rect 200 2165 215 2185
rect 235 2165 265 2185
rect 285 2165 300 2185
rect 200 2150 300 2165
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4585 600 4615
rect 550 4565 565 4585
rect 585 4565 600 4585
rect 550 4535 600 4565
rect 550 4515 565 4535
rect 585 4515 600 4535
rect 550 4485 600 4515
rect 550 4465 565 4485
rect 585 4465 600 4485
rect 550 4435 600 4465
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4335 600 4365
rect 550 4315 565 4335
rect 585 4315 600 4335
rect 550 4285 600 4315
rect 550 4265 565 4285
rect 585 4265 600 4285
rect 550 4235 600 4265
rect 550 4215 565 4235
rect 585 4215 600 4235
rect 550 4185 600 4215
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3935 600 3965
rect 550 3915 565 3935
rect 585 3915 600 3935
rect 550 3885 600 3915
rect 550 3865 565 3885
rect 585 3865 600 3885
rect 550 3835 600 3865
rect 550 3815 565 3835
rect 585 3815 600 3835
rect 550 3785 600 3815
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3685 600 3715
rect 550 3665 565 3685
rect 585 3665 600 3685
rect 550 3635 600 3665
rect 550 3615 565 3635
rect 585 3615 600 3635
rect 550 3585 600 3615
rect 550 3565 565 3585
rect 585 3565 600 3585
rect 550 3535 600 3565
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3285 600 3315
rect 550 3265 565 3285
rect 585 3265 600 3285
rect 550 3235 600 3265
rect 550 3215 565 3235
rect 585 3215 600 3235
rect 550 3185 600 3215
rect 550 3165 565 3185
rect 585 3165 600 3185
rect 550 3135 600 3165
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3035 600 3065
rect 550 3015 565 3035
rect 585 3015 600 3035
rect 550 2985 600 3015
rect 550 2965 565 2985
rect 585 2965 600 2985
rect 550 2935 600 2965
rect 550 2915 565 2935
rect 585 2915 600 2935
rect 550 2885 600 2915
rect 550 2865 565 2885
rect 585 2865 600 2885
rect 550 2835 600 2865
rect 550 2815 565 2835
rect 585 2815 600 2835
rect 550 2785 600 2815
rect 550 2765 565 2785
rect 585 2765 600 2785
rect 550 2735 600 2765
rect 550 2715 565 2735
rect 585 2715 600 2735
rect 550 2685 600 2715
rect 550 2665 565 2685
rect 585 2665 600 2685
rect 550 2635 600 2665
rect 550 2615 565 2635
rect 585 2615 600 2635
rect 550 2585 600 2615
rect 550 2565 565 2585
rect 585 2565 600 2585
rect 550 2535 600 2565
rect 550 2515 565 2535
rect 585 2515 600 2535
rect 550 2485 600 2515
rect 550 2465 565 2485
rect 585 2465 600 2485
rect 550 2435 600 2465
rect 550 2415 565 2435
rect 585 2415 600 2435
rect 550 2385 600 2415
rect 550 2365 565 2385
rect 585 2365 600 2385
rect 550 2335 600 2365
rect 550 2315 565 2335
rect 585 2315 600 2335
rect 550 2285 600 2315
rect 550 2265 565 2285
rect 585 2265 600 2285
rect 550 2235 600 2265
rect 550 2215 565 2235
rect 585 2215 600 2235
rect 550 2185 600 2215
rect 550 2165 565 2185
rect 585 2165 600 2185
rect 550 2135 600 2165
rect 550 2115 565 2135
rect 585 2115 600 2135
rect 550 2085 600 2115
rect 550 2065 565 2085
rect 585 2065 600 2085
rect 550 2035 600 2065
rect 550 2015 565 2035
rect 585 2015 600 2035
rect 550 1985 600 2015
rect 550 1965 565 1985
rect 585 1965 600 1985
rect 550 1935 600 1965
rect 550 1915 565 1935
rect 585 1915 600 1935
rect 550 1885 600 1915
rect 550 1865 565 1885
rect 585 1865 600 1885
rect 550 1835 600 1865
rect 550 1815 565 1835
rect 585 1815 600 1835
rect 550 1785 600 1815
rect 550 1765 565 1785
rect 585 1765 600 1785
rect 550 1735 600 1765
rect 550 1715 565 1735
rect 585 1715 600 1735
rect 550 1685 600 1715
rect 550 1665 565 1685
rect 585 1665 600 1685
rect 550 1635 600 1665
rect 550 1615 565 1635
rect 585 1615 600 1635
rect 550 1585 600 1615
rect 550 1565 565 1585
rect 585 1565 600 1585
rect 550 1535 600 1565
rect 550 1515 565 1535
rect 585 1515 600 1535
rect 550 1485 600 1515
rect 550 1465 565 1485
rect 585 1465 600 1485
rect 550 1435 600 1465
rect 550 1415 565 1435
rect 585 1415 600 1435
rect 550 1385 600 1415
rect 550 1365 565 1385
rect 585 1365 600 1385
rect 550 1335 600 1365
rect 550 1315 565 1335
rect 585 1315 600 1335
rect 550 1285 600 1315
rect 550 1265 565 1285
rect 585 1265 600 1285
rect 550 1235 600 1265
rect 550 1215 565 1235
rect 585 1215 600 1235
rect 550 1185 600 1215
rect 550 1165 565 1185
rect 585 1165 600 1185
rect 550 1150 600 1165
rect 200 1135 600 1150
rect 200 1115 215 1135
rect 235 1115 265 1135
rect 285 1115 315 1135
rect 335 1115 365 1135
rect 385 1115 415 1135
rect 435 1115 465 1135
rect 485 1115 515 1135
rect 535 1115 565 1135
rect 585 1115 600 1135
rect 200 1100 600 1115
<< nsubdiff >>
rect 200 4785 450 4800
rect 200 4765 215 4785
rect 235 4765 265 4785
rect 285 4765 315 4785
rect 335 4765 365 4785
rect 385 4765 415 4785
rect 435 4765 450 4785
rect 200 4750 450 4765
rect 400 4735 450 4750
rect 400 4715 415 4735
rect 435 4715 450 4735
rect 400 4685 450 4715
rect 400 4665 415 4685
rect 435 4665 450 4685
rect 400 4635 450 4665
rect 400 4615 415 4635
rect 435 4615 450 4635
rect 400 4585 450 4615
rect 400 4565 415 4585
rect 435 4565 450 4585
rect 400 4535 450 4565
rect 400 4515 415 4535
rect 435 4515 450 4535
rect 400 4485 450 4515
rect 400 4465 415 4485
rect 435 4465 450 4485
rect 400 4435 450 4465
rect 400 4415 415 4435
rect 435 4415 450 4435
rect 400 4385 450 4415
rect 400 4365 415 4385
rect 435 4365 450 4385
rect 400 4335 450 4365
rect 400 4315 415 4335
rect 435 4315 450 4335
rect 400 4285 450 4315
rect 400 4265 415 4285
rect 435 4265 450 4285
rect 400 4235 450 4265
rect 400 4215 415 4235
rect 435 4215 450 4235
rect 400 4185 450 4215
rect 400 4165 415 4185
rect 435 4165 450 4185
rect 400 4135 450 4165
rect 400 4115 415 4135
rect 435 4115 450 4135
rect 400 4085 450 4115
rect 400 4065 415 4085
rect 435 4065 450 4085
rect 400 4050 450 4065
rect 200 4035 450 4050
rect 200 4015 215 4035
rect 235 4015 265 4035
rect 285 4015 315 4035
rect 335 4015 365 4035
rect 385 4015 415 4035
rect 435 4015 450 4035
rect 200 4000 450 4015
rect 400 3985 450 4000
rect 400 3965 415 3985
rect 435 3965 450 3985
rect 400 3935 450 3965
rect 400 3915 415 3935
rect 435 3915 450 3935
rect 400 3885 450 3915
rect 400 3865 415 3885
rect 435 3865 450 3885
rect 400 3835 450 3865
rect 400 3815 415 3835
rect 435 3815 450 3835
rect 400 3785 450 3815
rect 400 3765 415 3785
rect 435 3765 450 3785
rect 400 3735 450 3765
rect 400 3715 415 3735
rect 435 3715 450 3735
rect 400 3685 450 3715
rect 400 3665 415 3685
rect 435 3665 450 3685
rect 400 3635 450 3665
rect 400 3615 415 3635
rect 435 3615 450 3635
rect 400 3585 450 3615
rect 400 3565 415 3585
rect 435 3565 450 3585
rect 400 3535 450 3565
rect 400 3515 415 3535
rect 435 3515 450 3535
rect 400 3485 450 3515
rect 400 3465 415 3485
rect 435 3465 450 3485
rect 400 3435 450 3465
rect 400 3415 415 3435
rect 435 3415 450 3435
rect 400 3385 450 3415
rect 400 3365 415 3385
rect 435 3365 450 3385
rect 400 3335 450 3365
rect 400 3315 415 3335
rect 435 3315 450 3335
rect 400 3285 450 3315
rect 400 3265 415 3285
rect 435 3265 450 3285
rect 400 3235 450 3265
rect 400 3215 415 3235
rect 435 3215 450 3235
rect 400 3185 450 3215
rect 400 3165 415 3185
rect 435 3165 450 3185
rect 400 3135 450 3165
rect 400 3115 415 3135
rect 435 3115 450 3135
rect 400 3085 450 3115
rect 400 3065 415 3085
rect 435 3065 450 3085
rect 400 3035 450 3065
rect 400 3015 415 3035
rect 435 3015 450 3035
rect 400 2985 450 3015
rect 400 2965 415 2985
rect 435 2965 450 2985
rect 400 2935 450 2965
rect 400 2915 415 2935
rect 435 2915 450 2935
rect 400 2885 450 2915
rect 400 2865 415 2885
rect 435 2865 450 2885
rect 400 2835 450 2865
rect 400 2815 415 2835
rect 435 2815 450 2835
rect 400 2785 450 2815
rect 400 2765 415 2785
rect 435 2765 450 2785
rect 400 2735 450 2765
rect 400 2715 415 2735
rect 435 2715 450 2735
rect 400 2685 450 2715
rect 400 2665 415 2685
rect 435 2665 450 2685
rect 400 2635 450 2665
rect 400 2615 415 2635
rect 435 2615 450 2635
rect 400 2585 450 2615
rect 400 2565 415 2585
rect 435 2565 450 2585
rect 400 2535 450 2565
rect 400 2515 415 2535
rect 435 2515 450 2535
rect 400 2485 450 2515
rect 400 2465 415 2485
rect 435 2465 450 2485
rect 400 2435 450 2465
rect 400 2415 415 2435
rect 435 2415 450 2435
rect 400 2385 450 2415
rect 400 2365 415 2385
rect 435 2365 450 2385
rect 400 2335 450 2365
rect 400 2315 415 2335
rect 435 2315 450 2335
rect 400 2285 450 2315
rect 400 2265 415 2285
rect 435 2265 450 2285
rect 400 2235 450 2265
rect 400 2215 415 2235
rect 435 2215 450 2235
rect 400 2185 450 2215
rect 400 2165 415 2185
rect 435 2165 450 2185
rect 400 2135 450 2165
rect 400 2115 415 2135
rect 435 2115 450 2135
rect 400 2085 450 2115
rect 400 2065 415 2085
rect 435 2065 450 2085
rect 400 2050 450 2065
rect 200 2035 450 2050
rect 200 2015 215 2035
rect 235 2015 265 2035
rect 285 2015 315 2035
rect 335 2015 365 2035
rect 385 2015 415 2035
rect 435 2015 450 2035
rect 200 2000 450 2015
rect 400 1985 450 2000
rect 400 1965 415 1985
rect 435 1965 450 1985
rect 400 1935 450 1965
rect 400 1915 415 1935
rect 435 1915 450 1935
rect 400 1885 450 1915
rect 400 1865 415 1885
rect 435 1865 450 1885
rect 400 1835 450 1865
rect 400 1815 415 1835
rect 435 1815 450 1835
rect 400 1785 450 1815
rect 400 1765 415 1785
rect 435 1765 450 1785
rect 400 1735 450 1765
rect 400 1715 415 1735
rect 435 1715 450 1735
rect 400 1685 450 1715
rect 400 1665 415 1685
rect 435 1665 450 1685
rect 400 1635 450 1665
rect 400 1615 415 1635
rect 435 1615 450 1635
rect 400 1585 450 1615
rect 400 1565 415 1585
rect 435 1565 450 1585
rect 400 1535 450 1565
rect 400 1515 415 1535
rect 435 1515 450 1535
rect 400 1485 450 1515
rect 400 1465 415 1485
rect 435 1465 450 1485
rect 400 1435 450 1465
rect 400 1415 415 1435
rect 435 1415 450 1435
rect 400 1385 450 1415
rect 400 1365 415 1385
rect 435 1365 450 1385
rect 400 1335 450 1365
rect 400 1315 415 1335
rect 435 1315 450 1335
rect 400 1300 450 1315
rect 200 1285 450 1300
rect 200 1265 215 1285
rect 235 1265 265 1285
rect 285 1265 315 1285
rect 335 1265 365 1285
rect 385 1265 415 1285
rect 435 1265 450 1285
rect 200 1250 450 1265
<< psubdiffcont >>
rect 215 4915 235 4935
rect 265 4915 285 4935
rect 315 4915 335 4935
rect 365 4915 385 4935
rect 415 4915 435 4935
rect 465 4915 485 4935
rect 515 4915 535 4935
rect 565 4915 585 4935
rect 565 4865 585 4885
rect 565 4815 585 4835
rect 215 3865 235 3885
rect 265 3865 285 3885
rect 265 3815 285 3835
rect 265 3765 285 3785
rect 265 3715 285 3735
rect 265 3665 285 3685
rect 265 3615 285 3635
rect 265 3565 285 3585
rect 265 3515 285 3535
rect 265 3465 285 3485
rect 265 3415 285 3435
rect 265 3365 285 3385
rect 265 3315 285 3335
rect 265 3265 285 3285
rect 265 3215 285 3235
rect 265 3165 285 3185
rect 265 3115 285 3135
rect 265 3065 285 3085
rect 265 3015 285 3035
rect 265 2965 285 2985
rect 265 2915 285 2935
rect 265 2865 285 2885
rect 265 2815 285 2835
rect 265 2765 285 2785
rect 265 2715 285 2735
rect 265 2665 285 2685
rect 265 2615 285 2635
rect 265 2565 285 2585
rect 265 2515 285 2535
rect 265 2465 285 2485
rect 265 2415 285 2435
rect 265 2365 285 2385
rect 265 2315 285 2335
rect 265 2265 285 2285
rect 265 2215 285 2235
rect 215 2165 235 2185
rect 265 2165 285 2185
rect 565 4765 585 4785
rect 565 4715 585 4735
rect 565 4665 585 4685
rect 565 4615 585 4635
rect 565 4565 585 4585
rect 565 4515 585 4535
rect 565 4465 585 4485
rect 565 4415 585 4435
rect 565 4365 585 4385
rect 565 4315 585 4335
rect 565 4265 585 4285
rect 565 4215 585 4235
rect 565 4165 585 4185
rect 565 4115 585 4135
rect 565 4065 585 4085
rect 565 4015 585 4035
rect 565 3965 585 3985
rect 565 3915 585 3935
rect 565 3865 585 3885
rect 565 3815 585 3835
rect 565 3765 585 3785
rect 565 3715 585 3735
rect 565 3665 585 3685
rect 565 3615 585 3635
rect 565 3565 585 3585
rect 565 3515 585 3535
rect 565 3465 585 3485
rect 565 3415 585 3435
rect 565 3365 585 3385
rect 565 3315 585 3335
rect 565 3265 585 3285
rect 565 3215 585 3235
rect 565 3165 585 3185
rect 565 3115 585 3135
rect 565 3065 585 3085
rect 565 3015 585 3035
rect 565 2965 585 2985
rect 565 2915 585 2935
rect 565 2865 585 2885
rect 565 2815 585 2835
rect 565 2765 585 2785
rect 565 2715 585 2735
rect 565 2665 585 2685
rect 565 2615 585 2635
rect 565 2565 585 2585
rect 565 2515 585 2535
rect 565 2465 585 2485
rect 565 2415 585 2435
rect 565 2365 585 2385
rect 565 2315 585 2335
rect 565 2265 585 2285
rect 565 2215 585 2235
rect 565 2165 585 2185
rect 565 2115 585 2135
rect 565 2065 585 2085
rect 565 2015 585 2035
rect 565 1965 585 1985
rect 565 1915 585 1935
rect 565 1865 585 1885
rect 565 1815 585 1835
rect 565 1765 585 1785
rect 565 1715 585 1735
rect 565 1665 585 1685
rect 565 1615 585 1635
rect 565 1565 585 1585
rect 565 1515 585 1535
rect 565 1465 585 1485
rect 565 1415 585 1435
rect 565 1365 585 1385
rect 565 1315 585 1335
rect 565 1265 585 1285
rect 565 1215 585 1235
rect 565 1165 585 1185
rect 215 1115 235 1135
rect 265 1115 285 1135
rect 315 1115 335 1135
rect 365 1115 385 1135
rect 415 1115 435 1135
rect 465 1115 485 1135
rect 515 1115 535 1135
rect 565 1115 585 1135
<< nsubdiffcont >>
rect 215 4765 235 4785
rect 265 4765 285 4785
rect 315 4765 335 4785
rect 365 4765 385 4785
rect 415 4765 435 4785
rect 415 4715 435 4735
rect 415 4665 435 4685
rect 415 4615 435 4635
rect 415 4565 435 4585
rect 415 4515 435 4535
rect 415 4465 435 4485
rect 415 4415 435 4435
rect 415 4365 435 4385
rect 415 4315 435 4335
rect 415 4265 435 4285
rect 415 4215 435 4235
rect 415 4165 435 4185
rect 415 4115 435 4135
rect 415 4065 435 4085
rect 215 4015 235 4035
rect 265 4015 285 4035
rect 315 4015 335 4035
rect 365 4015 385 4035
rect 415 4015 435 4035
rect 415 3965 435 3985
rect 415 3915 435 3935
rect 415 3865 435 3885
rect 415 3815 435 3835
rect 415 3765 435 3785
rect 415 3715 435 3735
rect 415 3665 435 3685
rect 415 3615 435 3635
rect 415 3565 435 3585
rect 415 3515 435 3535
rect 415 3465 435 3485
rect 415 3415 435 3435
rect 415 3365 435 3385
rect 415 3315 435 3335
rect 415 3265 435 3285
rect 415 3215 435 3235
rect 415 3165 435 3185
rect 415 3115 435 3135
rect 415 3065 435 3085
rect 415 3015 435 3035
rect 415 2965 435 2985
rect 415 2915 435 2935
rect 415 2865 435 2885
rect 415 2815 435 2835
rect 415 2765 435 2785
rect 415 2715 435 2735
rect 415 2665 435 2685
rect 415 2615 435 2635
rect 415 2565 435 2585
rect 415 2515 435 2535
rect 415 2465 435 2485
rect 415 2415 435 2435
rect 415 2365 435 2385
rect 415 2315 435 2335
rect 415 2265 435 2285
rect 415 2215 435 2235
rect 415 2165 435 2185
rect 415 2115 435 2135
rect 415 2065 435 2085
rect 215 2015 235 2035
rect 265 2015 285 2035
rect 315 2015 335 2035
rect 365 2015 385 2035
rect 415 2015 435 2035
rect 415 1965 435 1985
rect 415 1915 435 1935
rect 415 1865 435 1885
rect 415 1815 435 1835
rect 415 1765 435 1785
rect 415 1715 435 1735
rect 415 1665 435 1685
rect 415 1615 435 1635
rect 415 1565 435 1585
rect 415 1515 435 1535
rect 415 1465 435 1485
rect 415 1415 435 1435
rect 415 1365 435 1385
rect 415 1315 435 1335
rect 215 1265 235 1285
rect 265 1265 285 1285
rect 315 1265 335 1285
rect 365 1265 385 1285
rect 415 1265 435 1285
<< locali >>
rect 200 4935 600 4950
rect 200 4915 215 4935
rect 235 4915 265 4935
rect 285 4915 315 4935
rect 335 4915 365 4935
rect 385 4915 415 4935
rect 435 4915 465 4935
rect 485 4915 515 4935
rect 535 4915 565 4935
rect 585 4915 600 4935
rect 200 4900 600 4915
rect 550 4885 600 4900
rect 550 4865 565 4885
rect 585 4865 600 4885
rect 550 4835 600 4865
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 200 4785 450 4800
rect 200 4765 215 4785
rect 235 4765 265 4785
rect 285 4765 315 4785
rect 335 4765 365 4785
rect 385 4765 415 4785
rect 435 4765 450 4785
rect 200 4750 450 4765
rect 400 4735 450 4750
rect 400 4715 415 4735
rect 435 4715 450 4735
rect 400 4685 450 4715
rect 400 4665 415 4685
rect 435 4665 450 4685
rect 400 4635 450 4665
rect 400 4615 415 4635
rect 435 4615 450 4635
rect 400 4585 450 4615
rect 400 4565 415 4585
rect 435 4565 450 4585
rect 400 4535 450 4565
rect 400 4515 415 4535
rect 435 4515 450 4535
rect 400 4485 450 4515
rect 400 4465 415 4485
rect 435 4465 450 4485
rect 400 4435 450 4465
rect 400 4415 415 4435
rect 435 4415 450 4435
rect 400 4385 450 4415
rect 400 4365 415 4385
rect 435 4365 450 4385
rect 400 4335 450 4365
rect 400 4315 415 4335
rect 435 4315 450 4335
rect 400 4285 450 4315
rect 400 4265 415 4285
rect 435 4265 450 4285
rect 400 4235 450 4265
rect 400 4215 415 4235
rect 435 4215 450 4235
rect 400 4185 450 4215
rect 400 4165 415 4185
rect 435 4165 450 4185
rect 400 4135 450 4165
rect 400 4115 415 4135
rect 435 4115 450 4135
rect 400 4085 450 4115
rect 400 4065 415 4085
rect 435 4065 450 4085
rect 400 4050 450 4065
rect 200 4035 450 4050
rect 200 4015 215 4035
rect 235 4015 265 4035
rect 285 4015 315 4035
rect 335 4015 365 4035
rect 385 4015 415 4035
rect 435 4015 450 4035
rect 200 4000 450 4015
rect 400 3985 450 4000
rect 400 3965 415 3985
rect 435 3965 450 3985
rect 400 3935 450 3965
rect 400 3915 415 3935
rect 435 3915 450 3935
rect 200 3885 300 3900
rect 200 3865 215 3885
rect 235 3865 265 3885
rect 285 3865 300 3885
rect 200 3850 300 3865
rect 250 3835 300 3850
rect 250 3815 265 3835
rect 285 3815 300 3835
rect 250 3785 300 3815
rect 250 3765 265 3785
rect 285 3765 300 3785
rect 250 3735 300 3765
rect 250 3715 265 3735
rect 285 3715 300 3735
rect 250 3685 300 3715
rect 250 3665 265 3685
rect 285 3665 300 3685
rect 250 3635 300 3665
rect 250 3615 265 3635
rect 285 3615 300 3635
rect 250 3585 300 3615
rect 250 3565 265 3585
rect 285 3565 300 3585
rect 250 3535 300 3565
rect 250 3515 265 3535
rect 285 3515 300 3535
rect 250 3485 300 3515
rect 250 3465 265 3485
rect 285 3465 300 3485
rect 250 3435 300 3465
rect 250 3415 265 3435
rect 285 3415 300 3435
rect 250 3385 300 3415
rect 250 3365 265 3385
rect 285 3365 300 3385
rect 250 3335 300 3365
rect 250 3315 265 3335
rect 285 3315 300 3335
rect 250 3285 300 3315
rect 250 3265 265 3285
rect 285 3265 300 3285
rect 250 3235 300 3265
rect 250 3215 265 3235
rect 285 3215 300 3235
rect 250 3185 300 3215
rect 250 3165 265 3185
rect 285 3165 300 3185
rect 250 3135 300 3165
rect 250 3115 265 3135
rect 285 3115 300 3135
rect 250 3085 300 3115
rect 250 3065 265 3085
rect 285 3065 300 3085
rect 250 3035 300 3065
rect 250 3015 265 3035
rect 285 3015 300 3035
rect 250 2985 300 3015
rect 250 2965 265 2985
rect 285 2965 300 2985
rect 250 2935 300 2965
rect 250 2915 265 2935
rect 285 2915 300 2935
rect 250 2885 300 2915
rect 250 2865 265 2885
rect 285 2865 300 2885
rect 250 2835 300 2865
rect 250 2815 265 2835
rect 285 2815 300 2835
rect 250 2785 300 2815
rect 250 2765 265 2785
rect 285 2765 300 2785
rect 250 2735 300 2765
rect 250 2715 265 2735
rect 285 2715 300 2735
rect 250 2685 300 2715
rect 250 2665 265 2685
rect 285 2665 300 2685
rect 250 2635 300 2665
rect 250 2615 265 2635
rect 285 2615 300 2635
rect 250 2585 300 2615
rect 250 2565 265 2585
rect 285 2565 300 2585
rect 250 2535 300 2565
rect 250 2515 265 2535
rect 285 2515 300 2535
rect 250 2485 300 2515
rect 250 2465 265 2485
rect 285 2465 300 2485
rect 250 2435 300 2465
rect 250 2415 265 2435
rect 285 2415 300 2435
rect 250 2385 300 2415
rect 250 2365 265 2385
rect 285 2365 300 2385
rect 250 2335 300 2365
rect 250 2315 265 2335
rect 285 2315 300 2335
rect 250 2285 300 2315
rect 250 2265 265 2285
rect 285 2265 300 2285
rect 250 2235 300 2265
rect 250 2215 265 2235
rect 285 2215 300 2235
rect 250 2200 300 2215
rect 200 2185 300 2200
rect 200 2165 215 2185
rect 235 2165 265 2185
rect 285 2165 300 2185
rect 200 2150 300 2165
rect 400 3885 450 3915
rect 400 3865 415 3885
rect 435 3865 450 3885
rect 400 3835 450 3865
rect 400 3815 415 3835
rect 435 3815 450 3835
rect 400 3785 450 3815
rect 400 3765 415 3785
rect 435 3765 450 3785
rect 400 3735 450 3765
rect 400 3715 415 3735
rect 435 3715 450 3735
rect 400 3685 450 3715
rect 400 3665 415 3685
rect 435 3665 450 3685
rect 400 3635 450 3665
rect 400 3615 415 3635
rect 435 3615 450 3635
rect 400 3585 450 3615
rect 400 3565 415 3585
rect 435 3565 450 3585
rect 400 3535 450 3565
rect 400 3515 415 3535
rect 435 3515 450 3535
rect 400 3485 450 3515
rect 400 3465 415 3485
rect 435 3465 450 3485
rect 400 3435 450 3465
rect 400 3415 415 3435
rect 435 3415 450 3435
rect 400 3385 450 3415
rect 400 3365 415 3385
rect 435 3365 450 3385
rect 400 3335 450 3365
rect 400 3315 415 3335
rect 435 3315 450 3335
rect 400 3285 450 3315
rect 400 3265 415 3285
rect 435 3265 450 3285
rect 400 3235 450 3265
rect 400 3215 415 3235
rect 435 3215 450 3235
rect 400 3185 450 3215
rect 400 3165 415 3185
rect 435 3165 450 3185
rect 400 3135 450 3165
rect 400 3115 415 3135
rect 435 3115 450 3135
rect 400 3085 450 3115
rect 400 3065 415 3085
rect 435 3065 450 3085
rect 400 3035 450 3065
rect 400 3015 415 3035
rect 435 3015 450 3035
rect 400 2985 450 3015
rect 400 2965 415 2985
rect 435 2965 450 2985
rect 400 2935 450 2965
rect 400 2915 415 2935
rect 435 2915 450 2935
rect 400 2885 450 2915
rect 400 2865 415 2885
rect 435 2865 450 2885
rect 400 2835 450 2865
rect 400 2815 415 2835
rect 435 2815 450 2835
rect 400 2785 450 2815
rect 400 2765 415 2785
rect 435 2765 450 2785
rect 400 2735 450 2765
rect 400 2715 415 2735
rect 435 2715 450 2735
rect 400 2685 450 2715
rect 400 2665 415 2685
rect 435 2665 450 2685
rect 400 2635 450 2665
rect 400 2615 415 2635
rect 435 2615 450 2635
rect 400 2585 450 2615
rect 400 2565 415 2585
rect 435 2565 450 2585
rect 400 2535 450 2565
rect 400 2515 415 2535
rect 435 2515 450 2535
rect 400 2485 450 2515
rect 400 2465 415 2485
rect 435 2465 450 2485
rect 400 2435 450 2465
rect 400 2415 415 2435
rect 435 2415 450 2435
rect 400 2385 450 2415
rect 400 2365 415 2385
rect 435 2365 450 2385
rect 400 2335 450 2365
rect 400 2315 415 2335
rect 435 2315 450 2335
rect 400 2285 450 2315
rect 400 2265 415 2285
rect 435 2265 450 2285
rect 400 2235 450 2265
rect 400 2215 415 2235
rect 435 2215 450 2235
rect 400 2185 450 2215
rect 400 2165 415 2185
rect 435 2165 450 2185
rect 400 2135 450 2165
rect 400 2115 415 2135
rect 435 2115 450 2135
rect 400 2085 450 2115
rect 400 2065 415 2085
rect 435 2065 450 2085
rect 400 2050 450 2065
rect 200 2035 450 2050
rect 200 2015 215 2035
rect 235 2015 265 2035
rect 285 2015 315 2035
rect 335 2015 365 2035
rect 385 2015 415 2035
rect 435 2015 450 2035
rect 200 2000 450 2015
rect 400 1985 450 2000
rect 400 1965 415 1985
rect 435 1965 450 1985
rect 400 1935 450 1965
rect 400 1915 415 1935
rect 435 1915 450 1935
rect 400 1885 450 1915
rect 400 1865 415 1885
rect 435 1865 450 1885
rect 400 1835 450 1865
rect 400 1815 415 1835
rect 435 1815 450 1835
rect 400 1785 450 1815
rect 400 1765 415 1785
rect 435 1765 450 1785
rect 400 1735 450 1765
rect 400 1715 415 1735
rect 435 1715 450 1735
rect 400 1685 450 1715
rect 400 1665 415 1685
rect 435 1665 450 1685
rect 400 1635 450 1665
rect 400 1615 415 1635
rect 435 1615 450 1635
rect 400 1585 450 1615
rect 400 1565 415 1585
rect 435 1565 450 1585
rect 400 1535 450 1565
rect 400 1515 415 1535
rect 435 1515 450 1535
rect 400 1485 450 1515
rect 400 1465 415 1485
rect 435 1465 450 1485
rect 400 1435 450 1465
rect 400 1415 415 1435
rect 435 1415 450 1435
rect 400 1385 450 1415
rect 400 1365 415 1385
rect 435 1365 450 1385
rect 400 1335 450 1365
rect 400 1315 415 1335
rect 435 1315 450 1335
rect 400 1300 450 1315
rect 200 1285 450 1300
rect 200 1265 215 1285
rect 235 1265 265 1285
rect 285 1265 315 1285
rect 335 1265 365 1285
rect 385 1265 415 1285
rect 435 1265 450 1285
rect 200 1250 450 1265
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4585 600 4615
rect 550 4565 565 4585
rect 585 4565 600 4585
rect 550 4535 600 4565
rect 550 4515 565 4535
rect 585 4515 600 4535
rect 550 4485 600 4515
rect 550 4465 565 4485
rect 585 4465 600 4485
rect 550 4435 600 4465
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4335 600 4365
rect 550 4315 565 4335
rect 585 4315 600 4335
rect 550 4285 600 4315
rect 550 4265 565 4285
rect 585 4265 600 4285
rect 550 4235 600 4265
rect 550 4215 565 4235
rect 585 4215 600 4235
rect 550 4185 600 4215
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3935 600 3965
rect 550 3915 565 3935
rect 585 3915 600 3935
rect 550 3885 600 3915
rect 550 3865 565 3885
rect 585 3865 600 3885
rect 550 3835 600 3865
rect 550 3815 565 3835
rect 585 3815 600 3835
rect 550 3785 600 3815
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3685 600 3715
rect 550 3665 565 3685
rect 585 3665 600 3685
rect 550 3635 600 3665
rect 550 3615 565 3635
rect 585 3615 600 3635
rect 550 3585 600 3615
rect 550 3565 565 3585
rect 585 3565 600 3585
rect 550 3535 600 3565
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3285 600 3315
rect 550 3265 565 3285
rect 585 3265 600 3285
rect 550 3235 600 3265
rect 550 3215 565 3235
rect 585 3215 600 3235
rect 550 3185 600 3215
rect 550 3165 565 3185
rect 585 3165 600 3185
rect 550 3135 600 3165
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3035 600 3065
rect 550 3015 565 3035
rect 585 3015 600 3035
rect 550 2985 600 3015
rect 550 2965 565 2985
rect 585 2965 600 2985
rect 550 2935 600 2965
rect 550 2915 565 2935
rect 585 2915 600 2935
rect 550 2885 600 2915
rect 550 2865 565 2885
rect 585 2865 600 2885
rect 550 2835 600 2865
rect 550 2815 565 2835
rect 585 2815 600 2835
rect 550 2785 600 2815
rect 550 2765 565 2785
rect 585 2765 600 2785
rect 550 2735 600 2765
rect 550 2715 565 2735
rect 585 2715 600 2735
rect 550 2685 600 2715
rect 550 2665 565 2685
rect 585 2665 600 2685
rect 550 2635 600 2665
rect 550 2615 565 2635
rect 585 2615 600 2635
rect 550 2585 600 2615
rect 550 2565 565 2585
rect 585 2565 600 2585
rect 550 2535 600 2565
rect 550 2515 565 2535
rect 585 2515 600 2535
rect 550 2485 600 2515
rect 550 2465 565 2485
rect 585 2465 600 2485
rect 550 2435 600 2465
rect 550 2415 565 2435
rect 585 2415 600 2435
rect 550 2385 600 2415
rect 550 2365 565 2385
rect 585 2365 600 2385
rect 550 2335 600 2365
rect 550 2315 565 2335
rect 585 2315 600 2335
rect 550 2285 600 2315
rect 550 2265 565 2285
rect 585 2265 600 2285
rect 550 2235 600 2265
rect 550 2215 565 2235
rect 585 2215 600 2235
rect 550 2185 600 2215
rect 550 2165 565 2185
rect 585 2165 600 2185
rect 550 2135 600 2165
rect 550 2115 565 2135
rect 585 2115 600 2135
rect 550 2085 600 2115
rect 550 2065 565 2085
rect 585 2065 600 2085
rect 550 2035 600 2065
rect 550 2015 565 2035
rect 585 2015 600 2035
rect 550 1985 600 2015
rect 550 1965 565 1985
rect 585 1965 600 1985
rect 550 1935 600 1965
rect 550 1915 565 1935
rect 585 1915 600 1935
rect 550 1885 600 1915
rect 550 1865 565 1885
rect 585 1865 600 1885
rect 550 1835 600 1865
rect 550 1815 565 1835
rect 585 1815 600 1835
rect 550 1785 600 1815
rect 550 1765 565 1785
rect 585 1765 600 1785
rect 550 1735 600 1765
rect 550 1715 565 1735
rect 585 1715 600 1735
rect 550 1685 600 1715
rect 550 1665 565 1685
rect 585 1665 600 1685
rect 550 1635 600 1665
rect 550 1615 565 1635
rect 585 1615 600 1635
rect 550 1585 600 1615
rect 550 1565 565 1585
rect 585 1565 600 1585
rect 550 1535 600 1565
rect 550 1515 565 1535
rect 585 1515 600 1535
rect 550 1485 600 1515
rect 550 1465 565 1485
rect 585 1465 600 1485
rect 550 1435 600 1465
rect 550 1415 565 1435
rect 585 1415 600 1435
rect 550 1385 600 1415
rect 550 1365 565 1385
rect 585 1365 600 1385
rect 550 1335 600 1365
rect 550 1315 565 1335
rect 585 1315 600 1335
rect 550 1285 600 1315
rect 550 1265 565 1285
rect 585 1265 600 1285
rect 550 1235 600 1265
rect 550 1215 565 1235
rect 585 1215 600 1235
rect 550 1185 600 1215
rect 550 1165 565 1185
rect 585 1165 600 1185
rect 550 1150 600 1165
rect 200 1135 600 1150
rect 200 1115 215 1135
rect 235 1115 265 1135
rect 285 1115 315 1135
rect 335 1115 365 1135
rect 385 1115 415 1135
rect 435 1115 465 1135
rect 485 1115 515 1135
rect 535 1115 565 1135
rect 585 1115 600 1135
rect 200 1100 600 1115
<< metal2 >>
rect 200 4800 600 4850
rect 200 4700 600 4750
rect 200 4600 600 4650
rect 200 4500 600 4550
rect 200 4400 600 4450
rect 200 4300 600 4350
rect 200 4200 600 4250
rect 200 4000 600 4050
rect 200 3900 600 3950
rect 200 3500 600 3550
rect 200 3400 600 3450
rect 200 3300 600 3350
rect 200 3200 600 3250
rect 200 3100 600 3150
rect 200 2900 600 2950
rect 200 2800 600 2850
rect 200 2700 600 2750
rect 200 2600 600 2650
rect 200 2500 600 2550
rect 200 2100 600 2150
rect 200 2000 600 2050
rect 200 1800 600 1850
rect 200 1700 600 1750
rect 200 1600 600 1650
rect 200 1500 600 1550
rect 200 1400 600 1450
rect 200 1300 600 1350
rect 200 1200 600 1250
<< metal3 >>
rect 200 4800 600 4850
rect 200 4700 600 4750
rect 200 4600 600 4650
rect 200 4500 600 4550
rect 200 4400 600 4450
rect 200 4300 600 4350
rect 200 4200 600 4250
rect 200 4000 600 4050
rect 200 3900 600 3950
rect 200 3500 600 3550
rect 200 3300 600 3350
rect 200 3100 600 3150
rect 200 2900 600 2950
rect 200 2700 600 2750
rect 200 2500 600 2550
rect 200 2100 600 2150
rect 200 2000 600 2050
rect 200 1800 600 1850
rect 200 1700 600 1750
rect 200 1600 600 1650
rect 200 1500 600 1550
rect 200 1400 600 1450
rect 200 1300 600 1350
rect 200 1200 600 1250
<< end >>
