* NGSPICE file created from ddaa.ext - technology: sky130A

.subckt invdummy bp bn vdd vss vsub
X0 vdd xpb xpb bp sky130_fd_pr__pfet_01v8_lvt ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=0.5
X1 xpt xpt vdd bp sky130_fd_pr__pfet_01v8_lvt ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=0.5
X2 vdd xpt xpt bp sky130_fd_pr__pfet_01v8_lvt ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=0.5
X3 xn xn vss bn sky130_fd_pr__nfet_01v8_lvt ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=0.5
X4 xpb xpb vdd bp sky130_fd_pr__pfet_01v8_lvt ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=0.5
X5 vss xn xn bn sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=0.5
X6 xn xn vss bn sky130_fd_pr__nfet_01v8_lvt ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=0.5
X7 vss xn xn bn sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=0.5
.ends

.subckt inv1p1 in out bp bn vreg vss vsub
X0 vreg in out bp sky130_fd_pr__pfet_01v8_lvt ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=4
X1 out in vreg bp sky130_fd_pr__pfet_01v8_lvt ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=4
X2 out in xt bn sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=4
X3 out in xb bn sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=4
X4 out in vreg bp sky130_fd_pr__pfet_01v8_lvt ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=4
X5 xt in vss bn sky130_fd_pr__nfet_01v8 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=4
X6 vreg in out bp sky130_fd_pr__pfet_01v8_lvt ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=4
X7 xb in vss bn sky130_fd_pr__nfet_01v8 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=4
.ends

.subckt ddaa_slice im op vreg om bn ip SUB vss bp
Xa0 ip om bp bn vreg vss SUB inv1p1
Xa1 om om bp bn vreg vss SUB inv1p1
Xa2 op om bp bn vreg vss SUB inv1p1
Xa3 ip om bp bn vreg vss SUB inv1p1
Xa4 im op bp bn vreg vss SUB inv1p1
Xa5 om op bp bn vreg vss SUB inv1p1
Xa6 op op bp bn vreg vss SUB inv1p1
Xa7 im op bp bn vreg vss SUB inv1p1
.ends

.subckt ddaa ipa ima ipb imb op om bp bn vdd vss vsub
Xinvdummy_0 bp bn vdd vss vsub invdummy
Xinvdummy_1 bp bn vdd vss vsub invdummy
Xinvdummy_5 bp bn vdd vss vsub invdummy
Xinvdummy_6 bp bn vdd vss vsub invdummy
Xddaa_slice_0 ima op vdd om bn ipa vsub vss bp ddaa_slice
Xddaa_slice_1 imb op vdd om bn ipb vsub vss bp ddaa_slice
Xddaa_slice_2 ima op vdd om bn ipa vsub vss bp ddaa_slice
Xddaa_slice_3 ima op vdd om bn ipa vsub vss bp ddaa_slice
Xddaa_slice_4 imb op vdd om bn ipb vsub vss bp ddaa_slice
Xddaa_slice_5 imb op vdd om bn ipb vsub vss bp ddaa_slice
.ends

