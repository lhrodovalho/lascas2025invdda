magic
tech sky130A
timestamp 1725186481
<< viali >>
rect -385 5765 -365 5785
rect -235 5765 -215 5785
rect -535 3865 -515 3885
rect 10265 3865 10285 3885
rect -535 3815 -515 3835
rect 10260 3810 10290 3840
rect -385 1915 -365 1935
rect -235 1915 -215 1935
<< metal1 >>
rect -400 5790 -350 5800
rect -400 5760 -390 5790
rect -360 5760 -350 5790
rect -400 5750 -350 5760
rect -250 5790 -200 5800
rect -250 5760 -240 5790
rect -210 5760 -200 5790
rect -250 5750 -200 5760
rect -550 3890 -500 3900
rect -550 3860 -540 3890
rect -510 3860 -500 3890
rect -550 3840 -500 3860
rect -550 3810 -540 3840
rect -510 3810 -500 3840
rect -550 3800 -500 3810
rect 10250 3890 10300 3900
rect 10250 3860 10260 3890
rect 10290 3860 10300 3890
rect 10250 3840 10300 3860
rect 10250 3810 10260 3840
rect 10290 3810 10300 3840
rect 10250 3800 10300 3810
rect -400 1940 -350 1950
rect -400 1910 -390 1940
rect -360 1910 -350 1940
rect -400 1900 -350 1910
rect -250 1940 -200 1950
rect -250 1910 -240 1940
rect -210 1910 -200 1940
rect -250 1900 -200 1910
<< via1 >>
rect -390 5785 -360 5790
rect -390 5765 -385 5785
rect -385 5765 -365 5785
rect -365 5765 -360 5785
rect -390 5760 -360 5765
rect -240 5785 -210 5790
rect -240 5765 -235 5785
rect -235 5765 -215 5785
rect -215 5765 -210 5785
rect -240 5760 -210 5765
rect -540 3885 -510 3890
rect -540 3865 -535 3885
rect -535 3865 -515 3885
rect -515 3865 -510 3885
rect -540 3860 -510 3865
rect -540 3835 -510 3840
rect -540 3815 -535 3835
rect -535 3815 -515 3835
rect -515 3815 -510 3835
rect -540 3810 -510 3815
rect 10260 3885 10290 3890
rect 10260 3865 10265 3885
rect 10265 3865 10285 3885
rect 10285 3865 10290 3885
rect 10260 3860 10290 3865
rect 10260 3810 10290 3840
rect -390 1935 -360 1940
rect -390 1915 -385 1935
rect -385 1915 -365 1935
rect -365 1915 -360 1935
rect -390 1910 -360 1915
rect -240 1935 -210 1940
rect -240 1915 -235 1935
rect -235 1915 -215 1935
rect -215 1915 -210 1935
rect -240 1910 -210 1915
<< metal2 >>
rect -400 5790 -350 5800
rect -400 5760 -390 5790
rect -360 5760 -350 5790
rect -400 5750 -350 5760
rect -250 5790 -200 5800
rect -250 5760 -240 5790
rect -210 5760 -200 5790
rect -250 5750 -200 5760
rect -1850 3890 11600 3900
rect -1850 3860 -1840 3890
rect -1810 3860 -540 3890
rect -510 3860 10260 3890
rect 10290 3860 11560 3890
rect 11590 3860 11600 3890
rect -1850 3840 11600 3860
rect -1850 3810 -1840 3840
rect -1810 3810 -540 3840
rect -510 3810 10260 3840
rect 10290 3810 11560 3840
rect 11590 3810 11600 3840
rect -1850 3800 11600 3810
rect -400 1940 -350 1950
rect -400 1910 -390 1940
rect -360 1910 -350 1940
rect -400 1900 -350 1910
rect -250 1940 -200 1950
rect -250 1910 -240 1940
rect -210 1910 -200 1940
rect -250 1900 -200 1910
<< via2 >>
rect -390 5760 -360 5790
rect -240 5760 -210 5790
rect -1840 3860 -1810 3890
rect -540 3860 -510 3890
rect 10260 3860 10290 3890
rect 11560 3860 11590 3890
rect -1840 3810 -1810 3840
rect -540 3810 -510 3840
rect 10260 3810 10290 3840
rect 11560 3810 11590 3840
rect -390 1910 -360 1940
rect -240 1910 -210 1940
<< metal3 >>
rect 11650 7645 16950 7650
rect 11650 7605 16805 7645
rect 16845 7605 16905 7645
rect 16945 7605 16950 7645
rect -1750 7595 -550 7600
rect -1750 7555 -1745 7595
rect -1705 7555 -1695 7595
rect -1655 7555 -1645 7595
rect -1605 7555 -1595 7595
rect -1555 7555 -1545 7595
rect -1505 7555 -550 7595
rect -1750 7550 -550 7555
rect 10300 7595 11500 7600
rect 10300 7555 11255 7595
rect 11295 7555 11305 7595
rect 11345 7555 11355 7595
rect 11395 7555 11405 7595
rect 11445 7555 11455 7595
rect 11495 7555 11500 7595
rect 10300 7550 11500 7555
rect 11650 7595 16950 7605
rect 11650 7555 16805 7595
rect 16845 7555 16905 7595
rect 16945 7555 16950 7595
rect 11650 7545 16950 7555
rect 11650 7505 16805 7545
rect 16845 7505 16905 7545
rect 16945 7505 16950 7545
rect -1750 7495 -550 7500
rect -1750 7455 -1745 7495
rect -1705 7455 -1695 7495
rect -1655 7455 -1645 7495
rect -1605 7455 -1595 7495
rect -1555 7455 -1545 7495
rect -1505 7455 -550 7495
rect -1750 7450 -550 7455
rect 10300 7495 11500 7500
rect 10300 7455 11255 7495
rect 11295 7455 11305 7495
rect 11345 7455 11355 7495
rect 11395 7455 11405 7495
rect 11445 7455 11455 7495
rect 11495 7455 11500 7495
rect 10300 7450 11500 7455
rect 11650 7495 16950 7505
rect 11650 7455 16805 7495
rect 16845 7455 16905 7495
rect 16945 7455 16950 7495
rect 11650 7445 16950 7455
rect 11650 7405 16805 7445
rect 16845 7405 16905 7445
rect 16945 7405 16950 7445
rect -1750 7395 -550 7400
rect -1750 7355 -1745 7395
rect -1705 7355 -1695 7395
rect -1655 7355 -1645 7395
rect -1605 7355 -1595 7395
rect -1555 7355 -1545 7395
rect -1505 7355 -550 7395
rect -1750 7350 -550 7355
rect 10300 7395 11500 7400
rect 10300 7355 11255 7395
rect 11295 7355 11305 7395
rect 11345 7355 11355 7395
rect 11395 7355 11405 7395
rect 11445 7355 11455 7395
rect 11495 7355 11500 7395
rect 10300 7350 11500 7355
rect 11650 7395 16950 7405
rect 11650 7355 16805 7395
rect 16845 7355 16905 7395
rect 16945 7355 16950 7395
rect 11650 7345 16950 7355
rect 11650 7305 16805 7345
rect 16845 7305 16905 7345
rect 16945 7305 16950 7345
rect -1750 7295 -550 7300
rect -1750 7255 -1745 7295
rect -1705 7255 -1695 7295
rect -1655 7255 -1645 7295
rect -1605 7255 -1595 7295
rect -1555 7255 -1545 7295
rect -1505 7255 -550 7295
rect -1750 7250 -550 7255
rect 10300 7295 11500 7300
rect 10300 7255 11255 7295
rect 11295 7255 11305 7295
rect 11345 7255 11355 7295
rect 11395 7255 11405 7295
rect 11445 7255 11455 7295
rect 11495 7255 11500 7295
rect 10300 7250 11500 7255
rect 11650 7295 16950 7305
rect 11650 7255 16805 7295
rect 16845 7255 16905 7295
rect 16945 7255 16950 7295
rect 11650 7245 16950 7255
rect 11650 7205 16805 7245
rect 16845 7205 16905 7245
rect 16945 7205 16950 7245
rect -1750 7195 -550 7200
rect -1750 7155 -1745 7195
rect -1705 7155 -1695 7195
rect -1655 7155 -1645 7195
rect -1605 7155 -1595 7195
rect -1555 7155 -1545 7195
rect -1505 7155 -550 7195
rect -1750 7150 -550 7155
rect 10300 7195 11500 7200
rect 10300 7155 11255 7195
rect 11295 7155 11305 7195
rect 11345 7155 11355 7195
rect 11395 7155 11405 7195
rect 11445 7155 11455 7195
rect 11495 7155 11500 7195
rect 10300 7150 11500 7155
rect 11650 7195 16950 7205
rect 11650 7155 16805 7195
rect 16845 7155 16905 7195
rect 16945 7155 16950 7195
rect 11650 7145 16950 7155
rect 11650 7105 16805 7145
rect 16845 7105 16905 7145
rect 16945 7105 16950 7145
rect -1750 7095 -550 7100
rect -1750 7055 -1745 7095
rect -1705 7055 -1695 7095
rect -1655 7055 -1645 7095
rect -1605 7055 -1595 7095
rect -1555 7055 -1545 7095
rect -1505 7055 -550 7095
rect -1750 7050 -550 7055
rect 10300 7095 11500 7100
rect 10300 7055 11255 7095
rect 11295 7055 11305 7095
rect 11345 7055 11355 7095
rect 11395 7055 11405 7095
rect 11445 7055 11455 7095
rect 11495 7055 11500 7095
rect 10300 7050 11500 7055
rect 11650 7095 16950 7105
rect 11650 7055 16805 7095
rect 16845 7055 16905 7095
rect 16945 7055 16950 7095
rect 11650 7045 16950 7055
rect 11650 7005 16805 7045
rect 16845 7005 16905 7045
rect 16945 7005 16950 7045
rect -1750 6995 -550 7000
rect -1750 6955 -1745 6995
rect -1705 6955 -1695 6995
rect -1655 6955 -1645 6995
rect -1605 6955 -1595 6995
rect -1555 6955 -1545 6995
rect -1505 6955 -550 6995
rect -1750 6950 -550 6955
rect 10300 6995 11500 7000
rect 10300 6955 11255 6995
rect 11295 6955 11305 6995
rect 11345 6955 11355 6995
rect 11395 6955 11405 6995
rect 11445 6955 11455 6995
rect 11495 6955 11500 6995
rect 10300 6950 11500 6955
rect 11650 6995 16950 7005
rect 11650 6955 16805 6995
rect 16845 6955 16905 6995
rect 16945 6955 16950 6995
rect 11650 6945 16950 6955
rect 11650 6905 16805 6945
rect 16845 6905 16905 6945
rect 16945 6905 16950 6945
rect 11650 6895 16950 6905
rect 11650 6855 16805 6895
rect 16845 6855 16905 6895
rect 16945 6855 16950 6895
rect 11650 6845 16950 6855
rect 11650 6805 16805 6845
rect 16845 6805 16905 6845
rect 16945 6805 16950 6845
rect 11650 6795 16950 6805
rect 11650 6755 16805 6795
rect 16845 6755 16905 6795
rect 16945 6755 16950 6795
rect 11650 6745 16950 6755
rect 11650 6705 16805 6745
rect 16845 6705 16905 6745
rect 16945 6705 16950 6745
rect -1450 6695 -550 6700
rect -1450 6655 -1445 6695
rect -1405 6655 -1245 6695
rect -1205 6655 -1045 6695
rect -1005 6655 -845 6695
rect -805 6655 -645 6695
rect -605 6655 -550 6695
rect -1450 6650 -550 6655
rect 10300 6695 11200 6700
rect 10300 6655 10355 6695
rect 10395 6655 10755 6695
rect 10795 6655 11155 6695
rect 11195 6655 11200 6695
rect 10300 6650 11200 6655
rect 11650 6695 16950 6705
rect 11650 6655 16805 6695
rect 16845 6655 16905 6695
rect 16945 6655 16950 6695
rect 11650 6650 16950 6655
rect 16800 6645 16950 6650
rect 16800 6605 16805 6645
rect 16845 6605 16905 6645
rect 16945 6605 16950 6645
rect 9700 6595 16750 6600
rect 9700 6555 10455 6595
rect 10495 6555 10655 6595
rect 10695 6555 11655 6595
rect 11695 6555 11705 6595
rect 11745 6555 11755 6595
rect 11795 6555 11805 6595
rect 11845 6555 11855 6595
rect 11895 6555 16605 6595
rect 16645 6555 16655 6595
rect 16695 6555 16705 6595
rect 16745 6555 16750 6595
rect 9700 6550 16750 6555
rect 16800 6595 16950 6605
rect 16800 6555 16805 6595
rect 16845 6555 16905 6595
rect 16945 6555 16950 6595
rect 16800 6550 16950 6555
rect 16900 6545 16950 6550
rect 16900 6505 16905 6545
rect 16945 6505 16950 6545
rect 16900 6500 16950 6505
rect 9700 6495 16950 6500
rect 9700 6455 10555 6495
rect 10595 6455 16905 6495
rect 16945 6455 16950 6495
rect 9700 6450 16950 6455
rect 16900 6445 16950 6450
rect 16900 6405 16905 6445
rect 16945 6405 16950 6445
rect 16900 6400 16950 6405
rect 9700 6395 16750 6400
rect 9700 6355 10455 6395
rect 10495 6355 10655 6395
rect 10695 6355 11655 6395
rect 11695 6355 11705 6395
rect 11745 6355 11755 6395
rect 11795 6355 11805 6395
rect 11845 6355 11855 6395
rect 11895 6355 16605 6395
rect 16645 6355 16655 6395
rect 16695 6355 16705 6395
rect 16745 6355 16750 6395
rect 9700 6350 16750 6355
rect 16800 6395 16950 6400
rect 16800 6355 16805 6395
rect 16845 6355 16905 6395
rect 16945 6355 16950 6395
rect 16800 6345 16950 6355
rect 16800 6305 16805 6345
rect 16845 6305 16905 6345
rect 16945 6305 16950 6345
rect 16800 6300 16950 6305
rect -1450 6295 -550 6300
rect -1450 6255 -1445 6295
rect -1405 6255 -1245 6295
rect -1205 6255 -1045 6295
rect -1005 6255 -845 6295
rect -805 6255 -645 6295
rect -605 6255 -550 6295
rect -1450 6250 -550 6255
rect 10300 6295 11200 6300
rect 10300 6255 10355 6295
rect 10395 6255 10755 6295
rect 10795 6255 11155 6295
rect 11195 6255 11200 6295
rect 10300 6250 11200 6255
rect 11650 6295 16950 6300
rect 11650 6255 16805 6295
rect 16845 6255 16905 6295
rect 16945 6255 16950 6295
rect 11650 6245 16950 6255
rect 11650 6205 16805 6245
rect 16845 6205 16905 6245
rect 16945 6205 16950 6245
rect -1350 6195 9700 6200
rect -1350 6155 -945 6195
rect -905 6155 9700 6195
rect -1350 6150 9700 6155
rect 11650 6195 16950 6205
rect 11650 6155 16805 6195
rect 16845 6155 16905 6195
rect 16945 6155 16950 6195
rect 11650 6145 16950 6155
rect 11650 6105 16805 6145
rect 16845 6105 16905 6145
rect 16945 6105 16950 6145
rect -1450 6095 -550 6100
rect -1450 6055 -1445 6095
rect -1405 6055 -1245 6095
rect -1205 6055 -1045 6095
rect -1005 6055 -845 6095
rect -805 6055 -645 6095
rect -605 6055 -550 6095
rect -1450 6050 -550 6055
rect 11650 6095 16950 6105
rect 11650 6055 16805 6095
rect 16845 6055 16905 6095
rect 16945 6055 16950 6095
rect 11650 6045 16950 6055
rect 11650 6005 16805 6045
rect 16845 6005 16905 6045
rect 16945 6005 16950 6045
rect -1350 5995 9700 6000
rect -1350 5955 -1345 5995
rect -1305 5955 9700 5995
rect -1350 5950 9700 5955
rect 11650 5945 16950 6005
rect 11650 5905 16805 5945
rect 16845 5905 16905 5945
rect 16945 5905 16950 5945
rect -1450 5895 -550 5900
rect -1450 5855 -1445 5895
rect -1405 5855 -1245 5895
rect -1205 5855 -1045 5895
rect -1005 5855 -845 5895
rect -805 5855 -645 5895
rect -605 5855 -550 5895
rect -1450 5850 -550 5855
rect 11650 5895 16950 5905
rect 11650 5855 16805 5895
rect 16845 5855 16905 5895
rect 16945 5855 16950 5895
rect 11650 5850 16950 5855
rect -400 5795 -350 5800
rect -400 5755 -395 5795
rect -355 5755 -350 5795
rect -400 5750 -350 5755
rect -250 5795 -200 5800
rect -250 5755 -245 5795
rect -205 5755 -200 5795
rect -250 5750 -200 5755
rect -1450 5695 -550 5700
rect -1450 5655 -1445 5695
rect -1405 5655 -1245 5695
rect -1205 5655 -1045 5695
rect -1005 5655 -845 5695
rect -805 5655 -645 5695
rect -605 5655 -550 5695
rect -1450 5650 -550 5655
rect 11650 5695 16950 5700
rect 11650 5655 16805 5695
rect 16845 5655 16905 5695
rect 16945 5655 16950 5695
rect 11650 5645 16950 5655
rect 11650 5605 16805 5645
rect 16845 5605 16905 5645
rect 16945 5605 16950 5645
rect -1350 5595 9700 5600
rect -1350 5555 -1145 5595
rect -1105 5555 9700 5595
rect -1350 5550 9700 5555
rect 11650 5545 16950 5605
rect 11650 5505 16805 5545
rect 16845 5505 16905 5545
rect 16945 5505 16950 5545
rect -1450 5495 -550 5500
rect -1450 5455 -1445 5495
rect -1405 5455 -1245 5495
rect -1205 5455 -1045 5495
rect -1005 5455 -845 5495
rect -805 5455 -645 5495
rect -605 5455 -550 5495
rect -1450 5450 -550 5455
rect 11650 5495 16950 5505
rect 11650 5455 16805 5495
rect 16845 5455 16905 5495
rect 16945 5455 16950 5495
rect 11650 5445 16950 5455
rect 11650 5405 16805 5445
rect 16845 5405 16905 5445
rect 16945 5405 16950 5445
rect -1350 5395 9700 5400
rect -1350 5355 -745 5395
rect -705 5355 9700 5395
rect -1350 5350 9700 5355
rect 11650 5395 16950 5405
rect 11650 5355 16805 5395
rect 16845 5355 16905 5395
rect 16945 5355 16950 5395
rect 11650 5345 16950 5355
rect 11650 5305 16805 5345
rect 16845 5305 16905 5345
rect 16945 5305 16950 5345
rect -1450 5295 -550 5300
rect -1450 5255 -1445 5295
rect -1405 5255 -1245 5295
rect -1205 5255 -1045 5295
rect -1005 5255 -845 5295
rect -805 5255 -645 5295
rect -605 5255 -550 5295
rect -1450 5250 -550 5255
rect 10300 5295 11200 5300
rect 10300 5255 10355 5295
rect 10395 5255 10755 5295
rect 10795 5255 11155 5295
rect 11195 5255 11200 5295
rect 10300 5250 11200 5255
rect 11650 5295 16950 5305
rect 11650 5255 16805 5295
rect 16845 5255 16905 5295
rect 16945 5255 16950 5295
rect 11650 5250 16950 5255
rect 16800 5245 16950 5250
rect 16800 5205 16805 5245
rect 16845 5205 16905 5245
rect 16945 5205 16950 5245
rect 9700 5195 16750 5200
rect 9700 5155 10855 5195
rect 10895 5155 11055 5195
rect 11095 5155 11655 5195
rect 11695 5155 11705 5195
rect 11745 5155 11755 5195
rect 11795 5155 11805 5195
rect 11845 5155 11855 5195
rect 11895 5155 16605 5195
rect 16645 5155 16655 5195
rect 16695 5155 16705 5195
rect 16745 5155 16750 5195
rect 9700 5150 16750 5155
rect 16800 5195 16950 5205
rect 16800 5155 16805 5195
rect 16845 5155 16905 5195
rect 16945 5155 16950 5195
rect 16800 5150 16950 5155
rect 16900 5145 16950 5150
rect 16900 5105 16905 5145
rect 16945 5105 16950 5145
rect 16900 5100 16950 5105
rect 9700 5095 16950 5100
rect 9700 5055 10955 5095
rect 10995 5055 16905 5095
rect 16945 5055 16950 5095
rect 9700 5050 16950 5055
rect 16900 5045 16950 5050
rect 16900 5005 16905 5045
rect 16945 5005 16950 5045
rect 16900 5000 16950 5005
rect 9700 4995 16750 5000
rect 9700 4955 10855 4995
rect 10895 4955 11055 4995
rect 11095 4955 11655 4995
rect 11695 4955 11705 4995
rect 11745 4955 11755 4995
rect 11795 4955 11805 4995
rect 11845 4955 11855 4995
rect 11895 4955 16605 4995
rect 16645 4955 16655 4995
rect 16695 4955 16705 4995
rect 16745 4955 16750 4995
rect 9700 4950 16750 4955
rect 16800 4995 16950 5000
rect 16800 4955 16805 4995
rect 16845 4955 16905 4995
rect 16945 4955 16950 4995
rect 16800 4945 16950 4955
rect 16800 4905 16805 4945
rect 16845 4905 16905 4945
rect 16945 4905 16950 4945
rect 16800 4900 16950 4905
rect -1450 4895 -550 4900
rect -1450 4855 -1445 4895
rect -1405 4855 -1245 4895
rect -1205 4855 -1045 4895
rect -1005 4855 -845 4895
rect -805 4855 -645 4895
rect -605 4855 -550 4895
rect -1450 4850 -550 4855
rect 10300 4895 11200 4900
rect 10300 4855 10355 4895
rect 10395 4855 10755 4895
rect 10795 4855 11155 4895
rect 11195 4855 11200 4895
rect 10300 4850 11200 4855
rect 11650 4895 16950 4900
rect 11650 4855 16805 4895
rect 16845 4855 16905 4895
rect 16945 4855 16950 4895
rect 11650 4845 16950 4855
rect 11650 4805 16805 4845
rect 16845 4805 16905 4845
rect 16945 4805 16950 4845
rect 11650 4795 16950 4805
rect 11650 4755 16805 4795
rect 16845 4755 16905 4795
rect 16945 4755 16950 4795
rect 11650 4745 16950 4755
rect 11650 4705 16805 4745
rect 16845 4705 16905 4745
rect 16945 4705 16950 4745
rect 11650 4695 16950 4705
rect 11650 4655 16805 4695
rect 16845 4655 16905 4695
rect 16945 4655 16950 4695
rect 11650 4645 16950 4655
rect 11650 4605 16805 4645
rect 16845 4605 16905 4645
rect 16945 4605 16950 4645
rect -1750 4595 -550 4600
rect -1750 4555 -1745 4595
rect -1705 4555 -1695 4595
rect -1655 4555 -1645 4595
rect -1605 4555 -1595 4595
rect -1555 4555 -1545 4595
rect -1505 4555 -550 4595
rect -1750 4550 -550 4555
rect 10300 4595 11500 4600
rect 10300 4555 11255 4595
rect 11295 4555 11305 4595
rect 11345 4555 11355 4595
rect 11395 4555 11405 4595
rect 11445 4555 11455 4595
rect 11495 4555 11500 4595
rect 10300 4550 11500 4555
rect 11650 4595 16950 4605
rect 11650 4555 16805 4595
rect 16845 4555 16905 4595
rect 16945 4555 16950 4595
rect 11650 4545 16950 4555
rect 11650 4505 16805 4545
rect 16845 4505 16905 4545
rect 16945 4505 16950 4545
rect -1750 4495 -550 4500
rect -1750 4455 -1745 4495
rect -1705 4455 -1695 4495
rect -1655 4455 -1645 4495
rect -1605 4455 -1595 4495
rect -1555 4455 -1545 4495
rect -1505 4455 -550 4495
rect -1750 4450 -550 4455
rect 10300 4495 11500 4500
rect 10300 4455 11255 4495
rect 11295 4455 11305 4495
rect 11345 4455 11355 4495
rect 11395 4455 11405 4495
rect 11445 4455 11455 4495
rect 11495 4455 11500 4495
rect 10300 4450 11500 4455
rect 11650 4495 16950 4505
rect 11650 4455 16805 4495
rect 16845 4455 16905 4495
rect 16945 4455 16950 4495
rect 11650 4445 16950 4455
rect 11650 4405 16805 4445
rect 16845 4405 16905 4445
rect 16945 4405 16950 4445
rect -1750 4395 -550 4400
rect -1750 4355 -1745 4395
rect -1705 4355 -1695 4395
rect -1655 4355 -1645 4395
rect -1605 4355 -1595 4395
rect -1555 4355 -1545 4395
rect -1505 4355 -550 4395
rect -1750 4350 -550 4355
rect 10300 4395 11500 4400
rect 10300 4355 11255 4395
rect 11295 4355 11305 4395
rect 11345 4355 11355 4395
rect 11395 4355 11405 4395
rect 11445 4355 11455 4395
rect 11495 4355 11500 4395
rect 10300 4350 11500 4355
rect 11650 4395 16950 4405
rect 11650 4355 16805 4395
rect 16845 4355 16905 4395
rect 16945 4355 16950 4395
rect 11650 4345 16950 4355
rect 11650 4305 16805 4345
rect 16845 4305 16905 4345
rect 16945 4305 16950 4345
rect -1750 4295 -550 4300
rect -1750 4255 -1745 4295
rect -1705 4255 -1695 4295
rect -1655 4255 -1645 4295
rect -1605 4255 -1595 4295
rect -1555 4255 -1545 4295
rect -1505 4255 -550 4295
rect -1750 4250 -550 4255
rect 10300 4295 11500 4300
rect 10300 4255 11255 4295
rect 11295 4255 11305 4295
rect 11345 4255 11355 4295
rect 11395 4255 11405 4295
rect 11445 4255 11455 4295
rect 11495 4255 11500 4295
rect 10300 4250 11500 4255
rect 11650 4295 16950 4305
rect 11650 4255 16805 4295
rect 16845 4255 16905 4295
rect 16945 4255 16950 4295
rect 11650 4245 16950 4255
rect 11650 4205 16805 4245
rect 16845 4205 16905 4245
rect 16945 4205 16950 4245
rect -1750 4195 -550 4200
rect -1750 4155 -1745 4195
rect -1705 4155 -1695 4195
rect -1655 4155 -1645 4195
rect -1605 4155 -1595 4195
rect -1555 4155 -1545 4195
rect -1505 4155 -550 4195
rect -1750 4150 -550 4155
rect 10300 4195 11500 4200
rect 10300 4155 11255 4195
rect 11295 4155 11305 4195
rect 11345 4155 11355 4195
rect 11395 4155 11405 4195
rect 11445 4155 11455 4195
rect 11495 4155 11500 4195
rect 10300 4150 11500 4155
rect 11650 4195 16950 4205
rect 11650 4155 16805 4195
rect 16845 4155 16905 4195
rect 16945 4155 16950 4195
rect 11650 4145 16950 4155
rect 11650 4105 16805 4145
rect 16845 4105 16905 4145
rect 16945 4105 16950 4145
rect -1750 4095 -550 4100
rect -1750 4055 -1745 4095
rect -1705 4055 -1695 4095
rect -1655 4055 -1645 4095
rect -1605 4055 -1595 4095
rect -1555 4055 -1545 4095
rect -1505 4055 -550 4095
rect -1750 4050 -550 4055
rect 10300 4095 11500 4100
rect 10300 4055 11255 4095
rect 11295 4055 11305 4095
rect 11345 4055 11355 4095
rect 11395 4055 11405 4095
rect 11445 4055 11455 4095
rect 11495 4055 11500 4095
rect 10300 4050 11500 4055
rect 11650 4095 16950 4105
rect 11650 4055 16805 4095
rect 16845 4055 16905 4095
rect 16945 4055 16950 4095
rect 11650 4045 16950 4055
rect 11650 4005 16805 4045
rect 16845 4005 16905 4045
rect 16945 4005 16950 4045
rect -1750 3995 -550 4000
rect -1750 3955 -1745 3995
rect -1705 3955 -1695 3995
rect -1655 3955 -1645 3995
rect -1605 3955 -1595 3995
rect -1555 3955 -1545 3995
rect -1505 3955 -550 3995
rect -1750 3950 -550 3955
rect 10300 3995 11500 4000
rect 10300 3955 11255 3995
rect 11295 3955 11305 3995
rect 11345 3955 11355 3995
rect 11395 3955 11405 3995
rect 11445 3955 11455 3995
rect 11495 3955 11500 3995
rect 10300 3950 11500 3955
rect 11650 3995 16950 4005
rect 11650 3955 16805 3995
rect 16845 3955 16905 3995
rect 16945 3955 16950 3995
rect 11650 3945 16950 3955
rect 11650 3905 16805 3945
rect 16845 3905 16905 3945
rect 16945 3905 16950 3945
rect 11650 3900 16950 3905
rect -1850 3895 11600 3900
rect -1850 3855 -1845 3895
rect -1805 3890 11555 3895
rect -1805 3860 -540 3890
rect -510 3860 10260 3890
rect 10290 3860 11555 3890
rect -1805 3855 11555 3860
rect 11595 3855 11600 3895
rect -1850 3845 11600 3855
rect -1850 3805 -1845 3845
rect -1805 3840 11555 3845
rect -1805 3810 -540 3840
rect -510 3810 10260 3840
rect 10290 3810 11555 3840
rect -1805 3805 11555 3810
rect 11595 3805 11600 3845
rect -1850 3800 11600 3805
rect 11650 3795 16950 3800
rect 11650 3755 16805 3795
rect 16845 3755 16905 3795
rect 16945 3755 16950 3795
rect -1750 3745 -550 3750
rect -1750 3705 -1745 3745
rect -1705 3705 -1695 3745
rect -1655 3705 -1645 3745
rect -1605 3705 -1595 3745
rect -1555 3705 -1545 3745
rect -1505 3705 -550 3745
rect -1750 3700 -550 3705
rect 10300 3745 11500 3750
rect 10300 3705 11255 3745
rect 11295 3705 11305 3745
rect 11345 3705 11355 3745
rect 11395 3705 11405 3745
rect 11445 3705 11455 3745
rect 11495 3705 11500 3745
rect 10300 3700 11500 3705
rect 11650 3745 16950 3755
rect 11650 3705 16805 3745
rect 16845 3705 16905 3745
rect 16945 3705 16950 3745
rect 11650 3695 16950 3705
rect 11650 3655 16805 3695
rect 16845 3655 16905 3695
rect 16945 3655 16950 3695
rect -1750 3645 -550 3650
rect -1750 3605 -1745 3645
rect -1705 3605 -1695 3645
rect -1655 3605 -1645 3645
rect -1605 3605 -1595 3645
rect -1555 3605 -1545 3645
rect -1505 3605 -550 3645
rect -1750 3600 -550 3605
rect 10300 3645 11500 3650
rect 10300 3605 11255 3645
rect 11295 3605 11305 3645
rect 11345 3605 11355 3645
rect 11395 3605 11405 3645
rect 11445 3605 11455 3645
rect 11495 3605 11500 3645
rect 10300 3600 11500 3605
rect 11650 3645 16950 3655
rect 11650 3605 16805 3645
rect 16845 3605 16905 3645
rect 16945 3605 16950 3645
rect 11650 3595 16950 3605
rect 11650 3555 16805 3595
rect 16845 3555 16905 3595
rect 16945 3555 16950 3595
rect -1750 3545 -550 3550
rect -1750 3505 -1745 3545
rect -1705 3505 -1695 3545
rect -1655 3505 -1645 3545
rect -1605 3505 -1595 3545
rect -1555 3505 -1545 3545
rect -1505 3505 -550 3545
rect -1750 3500 -550 3505
rect 10300 3545 11500 3550
rect 10300 3505 11255 3545
rect 11295 3505 11305 3545
rect 11345 3505 11355 3545
rect 11395 3505 11405 3545
rect 11445 3505 11455 3545
rect 11495 3505 11500 3545
rect 10300 3500 11500 3505
rect 11650 3545 16950 3555
rect 11650 3505 16805 3545
rect 16845 3505 16905 3545
rect 16945 3505 16950 3545
rect 11650 3495 16950 3505
rect 11650 3455 16805 3495
rect 16845 3455 16905 3495
rect 16945 3455 16950 3495
rect -1750 3445 -550 3450
rect -1750 3405 -1745 3445
rect -1705 3405 -1695 3445
rect -1655 3405 -1645 3445
rect -1605 3405 -1595 3445
rect -1555 3405 -1545 3445
rect -1505 3405 -550 3445
rect -1750 3400 -550 3405
rect 10300 3445 11500 3450
rect 10300 3405 11255 3445
rect 11295 3405 11305 3445
rect 11345 3405 11355 3445
rect 11395 3405 11405 3445
rect 11445 3405 11455 3445
rect 11495 3405 11500 3445
rect 10300 3400 11500 3405
rect 11650 3445 16950 3455
rect 11650 3405 16805 3445
rect 16845 3405 16905 3445
rect 16945 3405 16950 3445
rect 11650 3395 16950 3405
rect 11650 3355 16805 3395
rect 16845 3355 16905 3395
rect 16945 3355 16950 3395
rect -1750 3345 -550 3350
rect -1750 3305 -1745 3345
rect -1705 3305 -1695 3345
rect -1655 3305 -1645 3345
rect -1605 3305 -1595 3345
rect -1555 3305 -1545 3345
rect -1505 3305 -550 3345
rect -1750 3300 -550 3305
rect 10300 3345 11500 3350
rect 10300 3305 11255 3345
rect 11295 3305 11305 3345
rect 11345 3305 11355 3345
rect 11395 3305 11405 3345
rect 11445 3305 11455 3345
rect 11495 3305 11500 3345
rect 10300 3300 11500 3305
rect 11650 3345 16950 3355
rect 11650 3305 16805 3345
rect 16845 3305 16905 3345
rect 16945 3305 16950 3345
rect 11650 3295 16950 3305
rect 11650 3255 16805 3295
rect 16845 3255 16905 3295
rect 16945 3255 16950 3295
rect -1750 3245 -550 3250
rect -1750 3205 -1745 3245
rect -1705 3205 -1695 3245
rect -1655 3205 -1645 3245
rect -1605 3205 -1595 3245
rect -1555 3205 -1545 3245
rect -1505 3205 -550 3245
rect -1750 3200 -550 3205
rect 10300 3245 11500 3250
rect 10300 3205 11255 3245
rect 11295 3205 11305 3245
rect 11345 3205 11355 3245
rect 11395 3205 11405 3245
rect 11445 3205 11455 3245
rect 11495 3205 11500 3245
rect 10300 3200 11500 3205
rect 11650 3245 16950 3255
rect 11650 3205 16805 3245
rect 16845 3205 16905 3245
rect 16945 3205 16950 3245
rect 11650 3195 16950 3205
rect 11650 3155 16805 3195
rect 16845 3155 16905 3195
rect 16945 3155 16950 3195
rect -1750 3145 -550 3150
rect -1750 3105 -1745 3145
rect -1705 3105 -1695 3145
rect -1655 3105 -1645 3145
rect -1605 3105 -1595 3145
rect -1555 3105 -1545 3145
rect -1505 3105 -550 3145
rect -1750 3100 -550 3105
rect 10300 3145 11500 3150
rect 10300 3105 11255 3145
rect 11295 3105 11305 3145
rect 11345 3105 11355 3145
rect 11395 3105 11405 3145
rect 11445 3105 11455 3145
rect 11495 3105 11500 3145
rect 10300 3100 11500 3105
rect 11650 3145 16950 3155
rect 11650 3105 16805 3145
rect 16845 3105 16905 3145
rect 16945 3105 16950 3145
rect 11650 3095 16950 3105
rect 11650 3055 16805 3095
rect 16845 3055 16905 3095
rect 16945 3055 16950 3095
rect 11650 3045 16950 3055
rect 11650 3005 16805 3045
rect 16845 3005 16905 3045
rect 16945 3005 16950 3045
rect 11650 2995 16950 3005
rect 11650 2955 16805 2995
rect 16845 2955 16905 2995
rect 16945 2955 16950 2995
rect 11650 2945 16950 2955
rect 11650 2905 16805 2945
rect 16845 2905 16905 2945
rect 16945 2905 16950 2945
rect 11650 2895 16950 2905
rect 11650 2855 16805 2895
rect 16845 2855 16905 2895
rect 16945 2855 16950 2895
rect -1450 2845 -550 2850
rect -1450 2805 -1445 2845
rect -1405 2805 -1245 2845
rect -1205 2805 -1045 2845
rect -1005 2805 -845 2845
rect -805 2805 -645 2845
rect -605 2805 -550 2845
rect -1450 2800 -550 2805
rect 10300 2845 11200 2850
rect 10300 2805 10355 2845
rect 10395 2805 10755 2845
rect 10795 2805 11155 2845
rect 11195 2805 11200 2845
rect 10300 2800 11200 2805
rect 11650 2845 16950 2855
rect 11650 2805 16805 2845
rect 16845 2805 16905 2845
rect 16945 2805 16950 2845
rect 11650 2800 16950 2805
rect 16800 2795 16950 2800
rect 16800 2755 16805 2795
rect 16845 2755 16905 2795
rect 16945 2755 16950 2795
rect 9700 2745 16750 2750
rect 9700 2705 10855 2745
rect 10895 2705 11055 2745
rect 11095 2705 11655 2745
rect 11695 2705 11705 2745
rect 11745 2705 11755 2745
rect 11795 2705 11805 2745
rect 11845 2705 11855 2745
rect 11895 2705 16605 2745
rect 16645 2705 16655 2745
rect 16695 2705 16705 2745
rect 16745 2705 16750 2745
rect 9700 2700 16750 2705
rect 16800 2745 16950 2755
rect 16800 2705 16805 2745
rect 16845 2705 16905 2745
rect 16945 2705 16950 2745
rect 16800 2700 16950 2705
rect 16900 2695 16950 2700
rect 16900 2655 16905 2695
rect 16945 2655 16950 2695
rect 16900 2650 16950 2655
rect 9700 2645 16950 2650
rect 9700 2605 10955 2645
rect 10995 2605 16905 2645
rect 16945 2605 16950 2645
rect 9700 2600 16950 2605
rect 16900 2595 16950 2600
rect 16900 2555 16905 2595
rect 16945 2555 16950 2595
rect 16900 2550 16950 2555
rect 9700 2545 16750 2550
rect 9700 2505 10855 2545
rect 10895 2505 11055 2545
rect 11095 2505 11655 2545
rect 11695 2505 11705 2545
rect 11745 2505 11755 2545
rect 11795 2505 11805 2545
rect 11845 2505 11855 2545
rect 11895 2505 16605 2545
rect 16645 2505 16655 2545
rect 16695 2505 16705 2545
rect 16745 2505 16750 2545
rect 9700 2500 16750 2505
rect 16800 2545 16950 2550
rect 16800 2505 16805 2545
rect 16845 2505 16905 2545
rect 16945 2505 16950 2545
rect 16800 2495 16950 2505
rect 16800 2455 16805 2495
rect 16845 2455 16905 2495
rect 16945 2455 16950 2495
rect 16800 2450 16950 2455
rect -1450 2445 -550 2450
rect -1450 2405 -1445 2445
rect -1405 2405 -1245 2445
rect -1205 2405 -1045 2445
rect -1005 2405 -845 2445
rect -805 2405 -645 2445
rect -605 2405 -550 2445
rect -1450 2400 -550 2405
rect 10300 2445 11200 2450
rect 10300 2405 10355 2445
rect 10395 2405 10755 2445
rect 10795 2405 11155 2445
rect 11195 2405 11200 2445
rect 10300 2400 11200 2405
rect 11650 2445 16950 2450
rect 11650 2405 16805 2445
rect 16845 2405 16905 2445
rect 16945 2405 16950 2445
rect 11650 2395 16950 2405
rect 11650 2355 16805 2395
rect 16845 2355 16905 2395
rect 16945 2355 16950 2395
rect -1350 2345 9700 2350
rect -1350 2305 -745 2345
rect -705 2305 9700 2345
rect -1350 2300 9700 2305
rect 11650 2345 16950 2355
rect 11650 2305 16805 2345
rect 16845 2305 16905 2345
rect 16945 2305 16950 2345
rect 11650 2295 16950 2305
rect 11650 2255 16805 2295
rect 16845 2255 16905 2295
rect 16945 2255 16950 2295
rect -1450 2245 -550 2250
rect -1450 2205 -1445 2245
rect -1405 2205 -1245 2245
rect -1205 2205 -1045 2245
rect -1005 2205 -845 2245
rect -805 2205 -645 2245
rect -605 2205 -550 2245
rect -1450 2200 -550 2205
rect 11650 2245 16950 2255
rect 11650 2205 16805 2245
rect 16845 2205 16905 2245
rect 16945 2205 16950 2245
rect 11650 2195 16950 2205
rect 11650 2155 16805 2195
rect 16845 2155 16905 2195
rect 16945 2155 16950 2195
rect -1350 2145 9700 2150
rect -1350 2105 -1145 2145
rect -1105 2105 9700 2145
rect -1350 2100 9700 2105
rect 11650 2145 16950 2155
rect 11650 2105 16805 2145
rect 16845 2105 16905 2145
rect 16945 2105 16950 2145
rect 11650 2095 16950 2105
rect 11650 2055 16805 2095
rect 16845 2055 16905 2095
rect 16945 2055 16950 2095
rect -1450 2045 -550 2050
rect -1450 2005 -1445 2045
rect -1405 2005 -1245 2045
rect -1205 2005 -1045 2045
rect -1005 2005 -845 2045
rect -805 2005 -645 2045
rect -605 2005 -550 2045
rect -1450 2000 -550 2005
rect 11650 2045 16950 2055
rect 11650 2005 16805 2045
rect 16845 2005 16905 2045
rect 16945 2005 16950 2045
rect 11650 2000 16950 2005
rect -400 1945 -350 1950
rect -400 1905 -395 1945
rect -355 1905 -350 1945
rect -400 1900 -350 1905
rect -250 1945 -200 1950
rect -250 1905 -245 1945
rect -205 1905 -200 1945
rect -250 1900 -200 1905
rect -1450 1845 -550 1850
rect -1450 1805 -1445 1845
rect -1405 1805 -1245 1845
rect -1205 1805 -1045 1845
rect -1005 1805 -845 1845
rect -805 1805 -645 1845
rect -605 1805 -550 1845
rect -1450 1800 -550 1805
rect 11650 1845 16950 1850
rect 11650 1805 16805 1845
rect 16845 1805 16905 1845
rect 16945 1805 16950 1845
rect 11650 1795 16950 1805
rect 11650 1755 16805 1795
rect 16845 1755 16905 1795
rect 16945 1755 16950 1795
rect -1350 1745 9700 1750
rect -1350 1705 -1345 1745
rect -1305 1705 9700 1745
rect -1350 1700 9700 1705
rect 11650 1745 16950 1755
rect 11650 1705 16805 1745
rect 16845 1705 16905 1745
rect 16945 1705 16950 1745
rect 11650 1695 16950 1705
rect 11650 1655 16805 1695
rect 16845 1655 16905 1695
rect 16945 1655 16950 1695
rect -1450 1645 -550 1650
rect -1450 1605 -1445 1645
rect -1405 1605 -1245 1645
rect -1205 1605 -1045 1645
rect -1005 1605 -845 1645
rect -805 1605 -645 1645
rect -605 1605 -550 1645
rect -1450 1600 -550 1605
rect 11650 1645 16950 1655
rect 11650 1605 16805 1645
rect 16845 1605 16905 1645
rect 16945 1605 16950 1645
rect 11650 1595 16950 1605
rect 11650 1555 16805 1595
rect 16845 1555 16905 1595
rect 16945 1555 16950 1595
rect -1350 1545 9700 1550
rect -1350 1505 -945 1545
rect -905 1505 9700 1545
rect -1350 1500 9700 1505
rect 11650 1545 16950 1555
rect 11650 1505 16805 1545
rect 16845 1505 16905 1545
rect 16945 1505 16950 1545
rect 11650 1495 16950 1505
rect 11650 1455 16805 1495
rect 16845 1455 16905 1495
rect 16945 1455 16950 1495
rect -1450 1445 -550 1450
rect -1450 1405 -1445 1445
rect -1405 1405 -1245 1445
rect -1205 1405 -1045 1445
rect -1005 1405 -845 1445
rect -805 1405 -645 1445
rect -605 1405 -550 1445
rect -1450 1400 -550 1405
rect 10300 1445 11200 1450
rect 10300 1405 10355 1445
rect 10395 1405 10755 1445
rect 10795 1405 11155 1445
rect 11195 1405 11200 1445
rect 10300 1400 11200 1405
rect 11650 1445 16950 1455
rect 11650 1405 16805 1445
rect 16845 1405 16905 1445
rect 16945 1405 16950 1445
rect 11650 1400 16950 1405
rect 16800 1395 16950 1400
rect 16800 1355 16805 1395
rect 16845 1355 16905 1395
rect 16945 1355 16950 1395
rect 9700 1345 16750 1350
rect 9700 1305 10455 1345
rect 10495 1305 10655 1345
rect 10695 1305 11655 1345
rect 11695 1305 11705 1345
rect 11745 1305 11755 1345
rect 11795 1305 11805 1345
rect 11845 1305 11855 1345
rect 11895 1305 16605 1345
rect 16645 1305 16655 1345
rect 16695 1305 16705 1345
rect 16745 1305 16750 1345
rect 9700 1300 16750 1305
rect 16800 1345 16950 1355
rect 16800 1305 16805 1345
rect 16845 1305 16905 1345
rect 16945 1305 16950 1345
rect 16800 1300 16950 1305
rect 16900 1295 16950 1300
rect 16900 1255 16905 1295
rect 16945 1255 16950 1295
rect 16900 1250 16950 1255
rect 9700 1245 16950 1250
rect 9700 1205 10555 1245
rect 10595 1205 16905 1245
rect 16945 1205 16950 1245
rect 9700 1200 16950 1205
rect 16900 1195 16950 1200
rect 16900 1155 16905 1195
rect 16945 1155 16950 1195
rect 16900 1150 16950 1155
rect 9700 1145 16750 1150
rect 9700 1105 10455 1145
rect 10495 1105 10655 1145
rect 10695 1105 11655 1145
rect 11695 1105 11705 1145
rect 11745 1105 11755 1145
rect 11795 1105 11805 1145
rect 11845 1105 11855 1145
rect 11895 1105 16605 1145
rect 16645 1105 16655 1145
rect 16695 1105 16705 1145
rect 16745 1105 16750 1145
rect 9700 1100 16750 1105
rect 16800 1145 16950 1150
rect 16800 1105 16805 1145
rect 16845 1105 16905 1145
rect 16945 1105 16950 1145
rect 16800 1095 16950 1105
rect 16800 1055 16805 1095
rect 16845 1055 16905 1095
rect 16945 1055 16950 1095
rect 16800 1050 16950 1055
rect -1450 1045 -550 1050
rect -1450 1005 -1445 1045
rect -1405 1005 -1245 1045
rect -1205 1005 -1045 1045
rect -1005 1005 -845 1045
rect -805 1005 -645 1045
rect -605 1005 -550 1045
rect -1450 1000 -550 1005
rect 10300 1045 11200 1050
rect 10300 1005 10355 1045
rect 10395 1005 10755 1045
rect 10795 1005 11155 1045
rect 11195 1005 11200 1045
rect 10300 1000 11200 1005
rect 11650 1045 16950 1050
rect 11650 1005 16805 1045
rect 16845 1005 16905 1045
rect 16945 1005 16950 1045
rect 11650 995 16950 1005
rect 11650 955 16805 995
rect 16845 955 16905 995
rect 16945 955 16950 995
rect 11650 945 16950 955
rect 11650 905 16805 945
rect 16845 905 16905 945
rect 16945 905 16950 945
rect 11650 895 16950 905
rect 11650 855 16805 895
rect 16845 855 16905 895
rect 16945 855 16950 895
rect 11650 845 16950 855
rect 11650 805 16805 845
rect 16845 805 16905 845
rect 16945 805 16950 845
rect 11650 795 16950 805
rect 11650 755 16805 795
rect 16845 755 16905 795
rect 16945 755 16950 795
rect -1750 745 -550 750
rect -1750 705 -1745 745
rect -1705 705 -1695 745
rect -1655 705 -1645 745
rect -1605 705 -1595 745
rect -1555 705 -1545 745
rect -1505 705 -550 745
rect -1750 700 -550 705
rect 10300 745 11500 750
rect 10300 705 11255 745
rect 11295 705 11305 745
rect 11345 705 11355 745
rect 11395 705 11405 745
rect 11445 705 11455 745
rect 11495 705 11500 745
rect 10300 700 11500 705
rect 11650 745 16950 755
rect 11650 705 16805 745
rect 16845 705 16905 745
rect 16945 705 16950 745
rect 11650 695 16950 705
rect 11650 655 16805 695
rect 16845 655 16905 695
rect 16945 655 16950 695
rect -1750 645 -550 650
rect -1750 605 -1745 645
rect -1705 605 -1695 645
rect -1655 605 -1645 645
rect -1605 605 -1595 645
rect -1555 605 -1545 645
rect -1505 605 -550 645
rect -1750 600 -550 605
rect 10300 645 11500 650
rect 10300 605 11255 645
rect 11295 605 11305 645
rect 11345 605 11355 645
rect 11395 605 11405 645
rect 11445 605 11455 645
rect 11495 605 11500 645
rect 10300 600 11500 605
rect 11650 645 16950 655
rect 11650 605 16805 645
rect 16845 605 16905 645
rect 16945 605 16950 645
rect 11650 595 16950 605
rect 11650 555 16805 595
rect 16845 555 16905 595
rect 16945 555 16950 595
rect -1750 545 -550 550
rect -1750 505 -1745 545
rect -1705 505 -1695 545
rect -1655 505 -1645 545
rect -1605 505 -1595 545
rect -1555 505 -1545 545
rect -1505 505 -550 545
rect -1750 500 -550 505
rect 10300 545 11500 550
rect 10300 505 11255 545
rect 11295 505 11305 545
rect 11345 505 11355 545
rect 11395 505 11405 545
rect 11445 505 11455 545
rect 11495 505 11500 545
rect 10300 500 11500 505
rect 11650 545 16950 555
rect 11650 505 16805 545
rect 16845 505 16905 545
rect 16945 505 16950 545
rect 11650 495 16950 505
rect 11650 455 16805 495
rect 16845 455 16905 495
rect 16945 455 16950 495
rect -1750 445 -550 450
rect -1750 405 -1745 445
rect -1705 405 -1695 445
rect -1655 405 -1645 445
rect -1605 405 -1595 445
rect -1555 405 -1545 445
rect -1505 405 -550 445
rect -1750 400 -550 405
rect 10300 445 11500 450
rect 10300 405 11255 445
rect 11295 405 11305 445
rect 11345 405 11355 445
rect 11395 405 11405 445
rect 11445 405 11455 445
rect 11495 405 11500 445
rect 10300 400 11500 405
rect 11650 445 16950 455
rect 11650 405 16805 445
rect 16845 405 16905 445
rect 16945 405 16950 445
rect 11650 395 16950 405
rect 11650 355 16805 395
rect 16845 355 16905 395
rect 16945 355 16950 395
rect -1750 345 -550 350
rect -1750 305 -1745 345
rect -1705 305 -1695 345
rect -1655 305 -1645 345
rect -1605 305 -1595 345
rect -1555 305 -1545 345
rect -1505 305 -550 345
rect -1750 300 -550 305
rect 10300 345 11500 350
rect 10300 305 11255 345
rect 11295 305 11305 345
rect 11345 305 11355 345
rect 11395 305 11405 345
rect 11445 305 11455 345
rect 11495 305 11500 345
rect 10300 300 11500 305
rect 11650 345 16950 355
rect 11650 305 16805 345
rect 16845 305 16905 345
rect 16945 305 16950 345
rect 11650 295 16950 305
rect 11650 255 16805 295
rect 16845 255 16905 295
rect 16945 255 16950 295
rect -1750 245 -550 250
rect -1750 205 -1745 245
rect -1705 205 -1695 245
rect -1655 205 -1645 245
rect -1605 205 -1595 245
rect -1555 205 -1545 245
rect -1505 205 -550 245
rect -1750 200 -550 205
rect 10300 245 11500 250
rect 10300 205 11255 245
rect 11295 205 11305 245
rect 11345 205 11355 245
rect 11395 205 11405 245
rect 11445 205 11455 245
rect 11495 205 11500 245
rect 10300 200 11500 205
rect 11650 245 16950 255
rect 11650 205 16805 245
rect 16845 205 16905 245
rect 16945 205 16950 245
rect 11650 195 16950 205
rect 11650 155 16805 195
rect 16845 155 16905 195
rect 16945 155 16950 195
rect -1750 145 -550 150
rect -1750 105 -1745 145
rect -1705 105 -1695 145
rect -1655 105 -1645 145
rect -1605 105 -1595 145
rect -1555 105 -1545 145
rect -1505 105 -550 145
rect -1750 100 -550 105
rect 10300 145 11500 150
rect 10300 105 11255 145
rect 11295 105 11305 145
rect 11345 105 11355 145
rect 11395 105 11405 145
rect 11445 105 11455 145
rect 11495 105 11500 145
rect 10300 100 11500 105
rect 11650 145 16950 155
rect 11650 105 16805 145
rect 16845 105 16905 145
rect 16945 105 16950 145
rect 11650 95 16950 105
rect 11650 55 16805 95
rect 16845 55 16905 95
rect 16945 55 16950 95
rect 11650 50 16950 55
<< via3 >>
rect 16805 7605 16845 7645
rect 16905 7605 16945 7645
rect -1745 7555 -1705 7595
rect -1695 7555 -1655 7595
rect -1645 7555 -1605 7595
rect -1595 7555 -1555 7595
rect -1545 7555 -1505 7595
rect 11255 7555 11295 7595
rect 11305 7555 11345 7595
rect 11355 7555 11395 7595
rect 11405 7555 11445 7595
rect 11455 7555 11495 7595
rect 16805 7555 16845 7595
rect 16905 7555 16945 7595
rect 16805 7505 16845 7545
rect 16905 7505 16945 7545
rect -1745 7455 -1705 7495
rect -1695 7455 -1655 7495
rect -1645 7455 -1605 7495
rect -1595 7455 -1555 7495
rect -1545 7455 -1505 7495
rect 11255 7455 11295 7495
rect 11305 7455 11345 7495
rect 11355 7455 11395 7495
rect 11405 7455 11445 7495
rect 11455 7455 11495 7495
rect 16805 7455 16845 7495
rect 16905 7455 16945 7495
rect 16805 7405 16845 7445
rect 16905 7405 16945 7445
rect -1745 7355 -1705 7395
rect -1695 7355 -1655 7395
rect -1645 7355 -1605 7395
rect -1595 7355 -1555 7395
rect -1545 7355 -1505 7395
rect 11255 7355 11295 7395
rect 11305 7355 11345 7395
rect 11355 7355 11395 7395
rect 11405 7355 11445 7395
rect 11455 7355 11495 7395
rect 16805 7355 16845 7395
rect 16905 7355 16945 7395
rect 16805 7305 16845 7345
rect 16905 7305 16945 7345
rect -1745 7255 -1705 7295
rect -1695 7255 -1655 7295
rect -1645 7255 -1605 7295
rect -1595 7255 -1555 7295
rect -1545 7255 -1505 7295
rect 11255 7255 11295 7295
rect 11305 7255 11345 7295
rect 11355 7255 11395 7295
rect 11405 7255 11445 7295
rect 11455 7255 11495 7295
rect 16805 7255 16845 7295
rect 16905 7255 16945 7295
rect 16805 7205 16845 7245
rect 16905 7205 16945 7245
rect -1745 7155 -1705 7195
rect -1695 7155 -1655 7195
rect -1645 7155 -1605 7195
rect -1595 7155 -1555 7195
rect -1545 7155 -1505 7195
rect 11255 7155 11295 7195
rect 11305 7155 11345 7195
rect 11355 7155 11395 7195
rect 11405 7155 11445 7195
rect 11455 7155 11495 7195
rect 16805 7155 16845 7195
rect 16905 7155 16945 7195
rect 16805 7105 16845 7145
rect 16905 7105 16945 7145
rect -1745 7055 -1705 7095
rect -1695 7055 -1655 7095
rect -1645 7055 -1605 7095
rect -1595 7055 -1555 7095
rect -1545 7055 -1505 7095
rect 11255 7055 11295 7095
rect 11305 7055 11345 7095
rect 11355 7055 11395 7095
rect 11405 7055 11445 7095
rect 11455 7055 11495 7095
rect 16805 7055 16845 7095
rect 16905 7055 16945 7095
rect 16805 7005 16845 7045
rect 16905 7005 16945 7045
rect -1745 6955 -1705 6995
rect -1695 6955 -1655 6995
rect -1645 6955 -1605 6995
rect -1595 6955 -1555 6995
rect -1545 6955 -1505 6995
rect 11255 6955 11295 6995
rect 11305 6955 11345 6995
rect 11355 6955 11395 6995
rect 11405 6955 11445 6995
rect 11455 6955 11495 6995
rect 16805 6955 16845 6995
rect 16905 6955 16945 6995
rect 16805 6905 16845 6945
rect 16905 6905 16945 6945
rect 16805 6855 16845 6895
rect 16905 6855 16945 6895
rect 16805 6805 16845 6845
rect 16905 6805 16945 6845
rect 16805 6755 16845 6795
rect 16905 6755 16945 6795
rect 16805 6705 16845 6745
rect 16905 6705 16945 6745
rect -1445 6655 -1405 6695
rect -1245 6655 -1205 6695
rect -1045 6655 -1005 6695
rect -845 6655 -805 6695
rect -645 6655 -605 6695
rect 10355 6655 10395 6695
rect 10755 6655 10795 6695
rect 11155 6655 11195 6695
rect 16805 6655 16845 6695
rect 16905 6655 16945 6695
rect 16805 6605 16845 6645
rect 16905 6605 16945 6645
rect 10455 6555 10495 6595
rect 10655 6555 10695 6595
rect 11655 6555 11695 6595
rect 11705 6555 11745 6595
rect 11755 6555 11795 6595
rect 11805 6555 11845 6595
rect 11855 6555 11895 6595
rect 16605 6555 16645 6595
rect 16655 6555 16695 6595
rect 16705 6555 16745 6595
rect 16805 6555 16845 6595
rect 16905 6555 16945 6595
rect 16905 6505 16945 6545
rect 10555 6455 10595 6495
rect 16905 6455 16945 6495
rect 16905 6405 16945 6445
rect 10455 6355 10495 6395
rect 10655 6355 10695 6395
rect 11655 6355 11695 6395
rect 11705 6355 11745 6395
rect 11755 6355 11795 6395
rect 11805 6355 11845 6395
rect 11855 6355 11895 6395
rect 16605 6355 16645 6395
rect 16655 6355 16695 6395
rect 16705 6355 16745 6395
rect 16805 6355 16845 6395
rect 16905 6355 16945 6395
rect 16805 6305 16845 6345
rect 16905 6305 16945 6345
rect -1445 6255 -1405 6295
rect -1245 6255 -1205 6295
rect -1045 6255 -1005 6295
rect -845 6255 -805 6295
rect -645 6255 -605 6295
rect 10355 6255 10395 6295
rect 10755 6255 10795 6295
rect 11155 6255 11195 6295
rect 16805 6255 16845 6295
rect 16905 6255 16945 6295
rect 16805 6205 16845 6245
rect 16905 6205 16945 6245
rect -945 6155 -905 6195
rect 16805 6155 16845 6195
rect 16905 6155 16945 6195
rect 16805 6105 16845 6145
rect 16905 6105 16945 6145
rect -1445 6055 -1405 6095
rect -1245 6055 -1205 6095
rect -1045 6055 -1005 6095
rect -845 6055 -805 6095
rect -645 6055 -605 6095
rect 16805 6055 16845 6095
rect 16905 6055 16945 6095
rect 16805 6005 16845 6045
rect 16905 6005 16945 6045
rect -1345 5955 -1305 5995
rect 16805 5905 16845 5945
rect 16905 5905 16945 5945
rect -1445 5855 -1405 5895
rect -1245 5855 -1205 5895
rect -1045 5855 -1005 5895
rect -845 5855 -805 5895
rect -645 5855 -605 5895
rect 16805 5855 16845 5895
rect 16905 5855 16945 5895
rect -395 5790 -355 5795
rect -395 5760 -390 5790
rect -390 5760 -360 5790
rect -360 5760 -355 5790
rect -395 5755 -355 5760
rect -245 5790 -205 5795
rect -245 5760 -240 5790
rect -240 5760 -210 5790
rect -210 5760 -205 5790
rect -245 5755 -205 5760
rect -1445 5655 -1405 5695
rect -1245 5655 -1205 5695
rect -1045 5655 -1005 5695
rect -845 5655 -805 5695
rect -645 5655 -605 5695
rect 16805 5655 16845 5695
rect 16905 5655 16945 5695
rect 16805 5605 16845 5645
rect 16905 5605 16945 5645
rect -1145 5555 -1105 5595
rect 16805 5505 16845 5545
rect 16905 5505 16945 5545
rect -1445 5455 -1405 5495
rect -1245 5455 -1205 5495
rect -1045 5455 -1005 5495
rect -845 5455 -805 5495
rect -645 5455 -605 5495
rect 16805 5455 16845 5495
rect 16905 5455 16945 5495
rect 16805 5405 16845 5445
rect 16905 5405 16945 5445
rect -745 5355 -705 5395
rect 16805 5355 16845 5395
rect 16905 5355 16945 5395
rect 16805 5305 16845 5345
rect 16905 5305 16945 5345
rect -1445 5255 -1405 5295
rect -1245 5255 -1205 5295
rect -1045 5255 -1005 5295
rect -845 5255 -805 5295
rect -645 5255 -605 5295
rect 10355 5255 10395 5295
rect 10755 5255 10795 5295
rect 11155 5255 11195 5295
rect 16805 5255 16845 5295
rect 16905 5255 16945 5295
rect 16805 5205 16845 5245
rect 16905 5205 16945 5245
rect 10855 5155 10895 5195
rect 11055 5155 11095 5195
rect 11655 5155 11695 5195
rect 11705 5155 11745 5195
rect 11755 5155 11795 5195
rect 11805 5155 11845 5195
rect 11855 5155 11895 5195
rect 16605 5155 16645 5195
rect 16655 5155 16695 5195
rect 16705 5155 16745 5195
rect 16805 5155 16845 5195
rect 16905 5155 16945 5195
rect 16905 5105 16945 5145
rect 10955 5055 10995 5095
rect 16905 5055 16945 5095
rect 16905 5005 16945 5045
rect 10855 4955 10895 4995
rect 11055 4955 11095 4995
rect 11655 4955 11695 4995
rect 11705 4955 11745 4995
rect 11755 4955 11795 4995
rect 11805 4955 11845 4995
rect 11855 4955 11895 4995
rect 16605 4955 16645 4995
rect 16655 4955 16695 4995
rect 16705 4955 16745 4995
rect 16805 4955 16845 4995
rect 16905 4955 16945 4995
rect 16805 4905 16845 4945
rect 16905 4905 16945 4945
rect -1445 4855 -1405 4895
rect -1245 4855 -1205 4895
rect -1045 4855 -1005 4895
rect -845 4855 -805 4895
rect -645 4855 -605 4895
rect 10355 4855 10395 4895
rect 10755 4855 10795 4895
rect 11155 4855 11195 4895
rect 16805 4855 16845 4895
rect 16905 4855 16945 4895
rect 16805 4805 16845 4845
rect 16905 4805 16945 4845
rect 16805 4755 16845 4795
rect 16905 4755 16945 4795
rect 16805 4705 16845 4745
rect 16905 4705 16945 4745
rect 16805 4655 16845 4695
rect 16905 4655 16945 4695
rect 16805 4605 16845 4645
rect 16905 4605 16945 4645
rect -1745 4555 -1705 4595
rect -1695 4555 -1655 4595
rect -1645 4555 -1605 4595
rect -1595 4555 -1555 4595
rect -1545 4555 -1505 4595
rect 11255 4555 11295 4595
rect 11305 4555 11345 4595
rect 11355 4555 11395 4595
rect 11405 4555 11445 4595
rect 11455 4555 11495 4595
rect 16805 4555 16845 4595
rect 16905 4555 16945 4595
rect 16805 4505 16845 4545
rect 16905 4505 16945 4545
rect -1745 4455 -1705 4495
rect -1695 4455 -1655 4495
rect -1645 4455 -1605 4495
rect -1595 4455 -1555 4495
rect -1545 4455 -1505 4495
rect 11255 4455 11295 4495
rect 11305 4455 11345 4495
rect 11355 4455 11395 4495
rect 11405 4455 11445 4495
rect 11455 4455 11495 4495
rect 16805 4455 16845 4495
rect 16905 4455 16945 4495
rect 16805 4405 16845 4445
rect 16905 4405 16945 4445
rect -1745 4355 -1705 4395
rect -1695 4355 -1655 4395
rect -1645 4355 -1605 4395
rect -1595 4355 -1555 4395
rect -1545 4355 -1505 4395
rect 11255 4355 11295 4395
rect 11305 4355 11345 4395
rect 11355 4355 11395 4395
rect 11405 4355 11445 4395
rect 11455 4355 11495 4395
rect 16805 4355 16845 4395
rect 16905 4355 16945 4395
rect 16805 4305 16845 4345
rect 16905 4305 16945 4345
rect -1745 4255 -1705 4295
rect -1695 4255 -1655 4295
rect -1645 4255 -1605 4295
rect -1595 4255 -1555 4295
rect -1545 4255 -1505 4295
rect 11255 4255 11295 4295
rect 11305 4255 11345 4295
rect 11355 4255 11395 4295
rect 11405 4255 11445 4295
rect 11455 4255 11495 4295
rect 16805 4255 16845 4295
rect 16905 4255 16945 4295
rect 16805 4205 16845 4245
rect 16905 4205 16945 4245
rect -1745 4155 -1705 4195
rect -1695 4155 -1655 4195
rect -1645 4155 -1605 4195
rect -1595 4155 -1555 4195
rect -1545 4155 -1505 4195
rect 11255 4155 11295 4195
rect 11305 4155 11345 4195
rect 11355 4155 11395 4195
rect 11405 4155 11445 4195
rect 11455 4155 11495 4195
rect 16805 4155 16845 4195
rect 16905 4155 16945 4195
rect 16805 4105 16845 4145
rect 16905 4105 16945 4145
rect -1745 4055 -1705 4095
rect -1695 4055 -1655 4095
rect -1645 4055 -1605 4095
rect -1595 4055 -1555 4095
rect -1545 4055 -1505 4095
rect 11255 4055 11295 4095
rect 11305 4055 11345 4095
rect 11355 4055 11395 4095
rect 11405 4055 11445 4095
rect 11455 4055 11495 4095
rect 16805 4055 16845 4095
rect 16905 4055 16945 4095
rect 16805 4005 16845 4045
rect 16905 4005 16945 4045
rect -1745 3955 -1705 3995
rect -1695 3955 -1655 3995
rect -1645 3955 -1605 3995
rect -1595 3955 -1555 3995
rect -1545 3955 -1505 3995
rect 11255 3955 11295 3995
rect 11305 3955 11345 3995
rect 11355 3955 11395 3995
rect 11405 3955 11445 3995
rect 11455 3955 11495 3995
rect 16805 3955 16845 3995
rect 16905 3955 16945 3995
rect 16805 3905 16845 3945
rect 16905 3905 16945 3945
rect -1845 3890 -1805 3895
rect 11555 3890 11595 3895
rect -1845 3860 -1840 3890
rect -1840 3860 -1810 3890
rect -1810 3860 -1805 3890
rect 11555 3860 11560 3890
rect 11560 3860 11590 3890
rect 11590 3860 11595 3890
rect -1845 3855 -1805 3860
rect 11555 3855 11595 3860
rect -1845 3840 -1805 3845
rect 11555 3840 11595 3845
rect -1845 3810 -1840 3840
rect -1840 3810 -1810 3840
rect -1810 3810 -1805 3840
rect 11555 3810 11560 3840
rect 11560 3810 11590 3840
rect 11590 3810 11595 3840
rect -1845 3805 -1805 3810
rect 11555 3805 11595 3810
rect 16805 3755 16845 3795
rect 16905 3755 16945 3795
rect -1745 3705 -1705 3745
rect -1695 3705 -1655 3745
rect -1645 3705 -1605 3745
rect -1595 3705 -1555 3745
rect -1545 3705 -1505 3745
rect 11255 3705 11295 3745
rect 11305 3705 11345 3745
rect 11355 3705 11395 3745
rect 11405 3705 11445 3745
rect 11455 3705 11495 3745
rect 16805 3705 16845 3745
rect 16905 3705 16945 3745
rect 16805 3655 16845 3695
rect 16905 3655 16945 3695
rect -1745 3605 -1705 3645
rect -1695 3605 -1655 3645
rect -1645 3605 -1605 3645
rect -1595 3605 -1555 3645
rect -1545 3605 -1505 3645
rect 11255 3605 11295 3645
rect 11305 3605 11345 3645
rect 11355 3605 11395 3645
rect 11405 3605 11445 3645
rect 11455 3605 11495 3645
rect 16805 3605 16845 3645
rect 16905 3605 16945 3645
rect 16805 3555 16845 3595
rect 16905 3555 16945 3595
rect -1745 3505 -1705 3545
rect -1695 3505 -1655 3545
rect -1645 3505 -1605 3545
rect -1595 3505 -1555 3545
rect -1545 3505 -1505 3545
rect 11255 3505 11295 3545
rect 11305 3505 11345 3545
rect 11355 3505 11395 3545
rect 11405 3505 11445 3545
rect 11455 3505 11495 3545
rect 16805 3505 16845 3545
rect 16905 3505 16945 3545
rect 16805 3455 16845 3495
rect 16905 3455 16945 3495
rect -1745 3405 -1705 3445
rect -1695 3405 -1655 3445
rect -1645 3405 -1605 3445
rect -1595 3405 -1555 3445
rect -1545 3405 -1505 3445
rect 11255 3405 11295 3445
rect 11305 3405 11345 3445
rect 11355 3405 11395 3445
rect 11405 3405 11445 3445
rect 11455 3405 11495 3445
rect 16805 3405 16845 3445
rect 16905 3405 16945 3445
rect 16805 3355 16845 3395
rect 16905 3355 16945 3395
rect -1745 3305 -1705 3345
rect -1695 3305 -1655 3345
rect -1645 3305 -1605 3345
rect -1595 3305 -1555 3345
rect -1545 3305 -1505 3345
rect 11255 3305 11295 3345
rect 11305 3305 11345 3345
rect 11355 3305 11395 3345
rect 11405 3305 11445 3345
rect 11455 3305 11495 3345
rect 16805 3305 16845 3345
rect 16905 3305 16945 3345
rect 16805 3255 16845 3295
rect 16905 3255 16945 3295
rect -1745 3205 -1705 3245
rect -1695 3205 -1655 3245
rect -1645 3205 -1605 3245
rect -1595 3205 -1555 3245
rect -1545 3205 -1505 3245
rect 11255 3205 11295 3245
rect 11305 3205 11345 3245
rect 11355 3205 11395 3245
rect 11405 3205 11445 3245
rect 11455 3205 11495 3245
rect 16805 3205 16845 3245
rect 16905 3205 16945 3245
rect 16805 3155 16845 3195
rect 16905 3155 16945 3195
rect -1745 3105 -1705 3145
rect -1695 3105 -1655 3145
rect -1645 3105 -1605 3145
rect -1595 3105 -1555 3145
rect -1545 3105 -1505 3145
rect 11255 3105 11295 3145
rect 11305 3105 11345 3145
rect 11355 3105 11395 3145
rect 11405 3105 11445 3145
rect 11455 3105 11495 3145
rect 16805 3105 16845 3145
rect 16905 3105 16945 3145
rect 16805 3055 16845 3095
rect 16905 3055 16945 3095
rect 16805 3005 16845 3045
rect 16905 3005 16945 3045
rect 16805 2955 16845 2995
rect 16905 2955 16945 2995
rect 16805 2905 16845 2945
rect 16905 2905 16945 2945
rect 16805 2855 16845 2895
rect 16905 2855 16945 2895
rect -1445 2805 -1405 2845
rect -1245 2805 -1205 2845
rect -1045 2805 -1005 2845
rect -845 2805 -805 2845
rect -645 2805 -605 2845
rect 10355 2805 10395 2845
rect 10755 2805 10795 2845
rect 11155 2805 11195 2845
rect 16805 2805 16845 2845
rect 16905 2805 16945 2845
rect 16805 2755 16845 2795
rect 16905 2755 16945 2795
rect 10855 2705 10895 2745
rect 11055 2705 11095 2745
rect 11655 2705 11695 2745
rect 11705 2705 11745 2745
rect 11755 2705 11795 2745
rect 11805 2705 11845 2745
rect 11855 2705 11895 2745
rect 16605 2705 16645 2745
rect 16655 2705 16695 2745
rect 16705 2705 16745 2745
rect 16805 2705 16845 2745
rect 16905 2705 16945 2745
rect 16905 2655 16945 2695
rect 10955 2605 10995 2645
rect 16905 2605 16945 2645
rect 16905 2555 16945 2595
rect 10855 2505 10895 2545
rect 11055 2505 11095 2545
rect 11655 2505 11695 2545
rect 11705 2505 11745 2545
rect 11755 2505 11795 2545
rect 11805 2505 11845 2545
rect 11855 2505 11895 2545
rect 16605 2505 16645 2545
rect 16655 2505 16695 2545
rect 16705 2505 16745 2545
rect 16805 2505 16845 2545
rect 16905 2505 16945 2545
rect 16805 2455 16845 2495
rect 16905 2455 16945 2495
rect -1445 2405 -1405 2445
rect -1245 2405 -1205 2445
rect -1045 2405 -1005 2445
rect -845 2405 -805 2445
rect -645 2405 -605 2445
rect 10355 2405 10395 2445
rect 10755 2405 10795 2445
rect 11155 2405 11195 2445
rect 16805 2405 16845 2445
rect 16905 2405 16945 2445
rect 16805 2355 16845 2395
rect 16905 2355 16945 2395
rect -745 2305 -705 2345
rect 16805 2305 16845 2345
rect 16905 2305 16945 2345
rect 16805 2255 16845 2295
rect 16905 2255 16945 2295
rect -1445 2205 -1405 2245
rect -1245 2205 -1205 2245
rect -1045 2205 -1005 2245
rect -845 2205 -805 2245
rect -645 2205 -605 2245
rect 16805 2205 16845 2245
rect 16905 2205 16945 2245
rect 16805 2155 16845 2195
rect 16905 2155 16945 2195
rect -1145 2105 -1105 2145
rect 16805 2105 16845 2145
rect 16905 2105 16945 2145
rect 16805 2055 16845 2095
rect 16905 2055 16945 2095
rect -1445 2005 -1405 2045
rect -1245 2005 -1205 2045
rect -1045 2005 -1005 2045
rect -845 2005 -805 2045
rect -645 2005 -605 2045
rect 16805 2005 16845 2045
rect 16905 2005 16945 2045
rect -395 1940 -355 1945
rect -395 1910 -390 1940
rect -390 1910 -360 1940
rect -360 1910 -355 1940
rect -395 1905 -355 1910
rect -245 1940 -205 1945
rect -245 1910 -240 1940
rect -240 1910 -210 1940
rect -210 1910 -205 1940
rect -245 1905 -205 1910
rect -1445 1805 -1405 1845
rect -1245 1805 -1205 1845
rect -1045 1805 -1005 1845
rect -845 1805 -805 1845
rect -645 1805 -605 1845
rect 16805 1805 16845 1845
rect 16905 1805 16945 1845
rect 16805 1755 16845 1795
rect 16905 1755 16945 1795
rect -1345 1705 -1305 1745
rect 16805 1705 16845 1745
rect 16905 1705 16945 1745
rect 16805 1655 16845 1695
rect 16905 1655 16945 1695
rect -1445 1605 -1405 1645
rect -1245 1605 -1205 1645
rect -1045 1605 -1005 1645
rect -845 1605 -805 1645
rect -645 1605 -605 1645
rect 16805 1605 16845 1645
rect 16905 1605 16945 1645
rect 16805 1555 16845 1595
rect 16905 1555 16945 1595
rect -945 1505 -905 1545
rect 16805 1505 16845 1545
rect 16905 1505 16945 1545
rect 16805 1455 16845 1495
rect 16905 1455 16945 1495
rect -1445 1405 -1405 1445
rect -1245 1405 -1205 1445
rect -1045 1405 -1005 1445
rect -845 1405 -805 1445
rect -645 1405 -605 1445
rect 10355 1405 10395 1445
rect 10755 1405 10795 1445
rect 11155 1405 11195 1445
rect 16805 1405 16845 1445
rect 16905 1405 16945 1445
rect 16805 1355 16845 1395
rect 16905 1355 16945 1395
rect 10455 1305 10495 1345
rect 10655 1305 10695 1345
rect 11655 1305 11695 1345
rect 11705 1305 11745 1345
rect 11755 1305 11795 1345
rect 11805 1305 11845 1345
rect 11855 1305 11895 1345
rect 16605 1305 16645 1345
rect 16655 1305 16695 1345
rect 16705 1305 16745 1345
rect 16805 1305 16845 1345
rect 16905 1305 16945 1345
rect 16905 1255 16945 1295
rect 10555 1205 10595 1245
rect 16905 1205 16945 1245
rect 16905 1155 16945 1195
rect 10455 1105 10495 1145
rect 10655 1105 10695 1145
rect 11655 1105 11695 1145
rect 11705 1105 11745 1145
rect 11755 1105 11795 1145
rect 11805 1105 11845 1145
rect 11855 1105 11895 1145
rect 16605 1105 16645 1145
rect 16655 1105 16695 1145
rect 16705 1105 16745 1145
rect 16805 1105 16845 1145
rect 16905 1105 16945 1145
rect 16805 1055 16845 1095
rect 16905 1055 16945 1095
rect -1445 1005 -1405 1045
rect -1245 1005 -1205 1045
rect -1045 1005 -1005 1045
rect -845 1005 -805 1045
rect -645 1005 -605 1045
rect 10355 1005 10395 1045
rect 10755 1005 10795 1045
rect 11155 1005 11195 1045
rect 16805 1005 16845 1045
rect 16905 1005 16945 1045
rect 16805 955 16845 995
rect 16905 955 16945 995
rect 16805 905 16845 945
rect 16905 905 16945 945
rect 16805 855 16845 895
rect 16905 855 16945 895
rect 16805 805 16845 845
rect 16905 805 16945 845
rect 16805 755 16845 795
rect 16905 755 16945 795
rect -1745 705 -1705 745
rect -1695 705 -1655 745
rect -1645 705 -1605 745
rect -1595 705 -1555 745
rect -1545 705 -1505 745
rect 11255 705 11295 745
rect 11305 705 11345 745
rect 11355 705 11395 745
rect 11405 705 11445 745
rect 11455 705 11495 745
rect 16805 705 16845 745
rect 16905 705 16945 745
rect 16805 655 16845 695
rect 16905 655 16945 695
rect -1745 605 -1705 645
rect -1695 605 -1655 645
rect -1645 605 -1605 645
rect -1595 605 -1555 645
rect -1545 605 -1505 645
rect 11255 605 11295 645
rect 11305 605 11345 645
rect 11355 605 11395 645
rect 11405 605 11445 645
rect 11455 605 11495 645
rect 16805 605 16845 645
rect 16905 605 16945 645
rect 16805 555 16845 595
rect 16905 555 16945 595
rect -1745 505 -1705 545
rect -1695 505 -1655 545
rect -1645 505 -1605 545
rect -1595 505 -1555 545
rect -1545 505 -1505 545
rect 11255 505 11295 545
rect 11305 505 11345 545
rect 11355 505 11395 545
rect 11405 505 11445 545
rect 11455 505 11495 545
rect 16805 505 16845 545
rect 16905 505 16945 545
rect 16805 455 16845 495
rect 16905 455 16945 495
rect -1745 405 -1705 445
rect -1695 405 -1655 445
rect -1645 405 -1605 445
rect -1595 405 -1555 445
rect -1545 405 -1505 445
rect 11255 405 11295 445
rect 11305 405 11345 445
rect 11355 405 11395 445
rect 11405 405 11445 445
rect 11455 405 11495 445
rect 16805 405 16845 445
rect 16905 405 16945 445
rect 16805 355 16845 395
rect 16905 355 16945 395
rect -1745 305 -1705 345
rect -1695 305 -1655 345
rect -1645 305 -1605 345
rect -1595 305 -1555 345
rect -1545 305 -1505 345
rect 11255 305 11295 345
rect 11305 305 11345 345
rect 11355 305 11395 345
rect 11405 305 11445 345
rect 11455 305 11495 345
rect 16805 305 16845 345
rect 16905 305 16945 345
rect 16805 255 16845 295
rect 16905 255 16945 295
rect -1745 205 -1705 245
rect -1695 205 -1655 245
rect -1645 205 -1605 245
rect -1595 205 -1555 245
rect -1545 205 -1505 245
rect 11255 205 11295 245
rect 11305 205 11345 245
rect 11355 205 11395 245
rect 11405 205 11445 245
rect 11455 205 11495 245
rect 16805 205 16845 245
rect 16905 205 16945 245
rect 16805 155 16845 195
rect 16905 155 16945 195
rect -1745 105 -1705 145
rect -1695 105 -1655 145
rect -1645 105 -1605 145
rect -1595 105 -1555 145
rect -1545 105 -1505 145
rect 11255 105 11295 145
rect 11305 105 11345 145
rect 11355 105 11395 145
rect 11405 105 11445 145
rect 11455 105 11495 145
rect 16805 105 16845 145
rect 16905 105 16945 145
rect 16805 55 16845 95
rect 16905 55 16945 95
<< mimcap >>
rect 11700 7550 16700 7600
rect 11700 6750 11750 7550
rect 16650 6750 16700 7550
rect 11700 6700 16700 6750
rect 11700 6200 16700 6250
rect 11700 5950 11750 6200
rect 16650 5950 16700 6200
rect 11700 5900 16700 5950
rect 11700 5600 16700 5650
rect 11700 5350 11750 5600
rect 16650 5350 16700 5600
rect 11700 5300 16700 5350
rect 11700 4800 16700 4850
rect 11700 4000 11750 4800
rect 16650 4000 16700 4800
rect 11700 3950 16700 4000
rect 11700 3700 16700 3750
rect 11700 2900 11750 3700
rect 16650 2900 16700 3700
rect 11700 2850 16700 2900
rect 11700 2350 16700 2400
rect 11700 2100 11750 2350
rect 16650 2100 16700 2350
rect 11700 2050 16700 2100
rect 11700 1750 16700 1800
rect 11700 1500 11750 1750
rect 16650 1500 16700 1750
rect 11700 1450 16700 1500
rect 11700 950 16700 1000
rect 11700 150 11750 950
rect 16650 150 16700 950
rect 11700 100 16700 150
<< mimcapcontact >>
rect 11750 6750 16650 7550
rect 11750 5950 16650 6200
rect 11750 5350 16650 5600
rect 11750 4000 16650 4800
rect 11750 2900 16650 3700
rect 11750 2100 16650 2350
rect 11750 1500 16650 1750
rect 11750 150 16650 950
<< metal4 >>
rect -1850 3895 -1800 7700
rect -1850 3855 -1845 3895
rect -1805 3855 -1800 3895
rect -1850 3845 -1800 3855
rect -1850 3805 -1845 3845
rect -1805 3805 -1800 3845
rect -1850 0 -1800 3805
rect -1750 7595 -1500 7700
rect -1750 7555 -1745 7595
rect -1705 7555 -1695 7595
rect -1655 7555 -1645 7595
rect -1605 7555 -1595 7595
rect -1555 7555 -1545 7595
rect -1505 7555 -1500 7595
rect -1750 7495 -1500 7555
rect -1750 7455 -1745 7495
rect -1705 7455 -1695 7495
rect -1655 7455 -1645 7495
rect -1605 7455 -1595 7495
rect -1555 7455 -1545 7495
rect -1505 7455 -1500 7495
rect -1750 7395 -1500 7455
rect -1750 7355 -1745 7395
rect -1705 7355 -1695 7395
rect -1655 7355 -1645 7395
rect -1605 7355 -1595 7395
rect -1555 7355 -1545 7395
rect -1505 7355 -1500 7395
rect -1750 7295 -1500 7355
rect -1750 7255 -1745 7295
rect -1705 7255 -1695 7295
rect -1655 7255 -1645 7295
rect -1605 7255 -1595 7295
rect -1555 7255 -1545 7295
rect -1505 7255 -1500 7295
rect -1750 7195 -1500 7255
rect -1750 7155 -1745 7195
rect -1705 7155 -1695 7195
rect -1655 7155 -1645 7195
rect -1605 7155 -1595 7195
rect -1555 7155 -1545 7195
rect -1505 7155 -1500 7195
rect -1750 7095 -1500 7155
rect -1750 7055 -1745 7095
rect -1705 7055 -1695 7095
rect -1655 7055 -1645 7095
rect -1605 7055 -1595 7095
rect -1555 7055 -1545 7095
rect -1505 7055 -1500 7095
rect -1750 6995 -1500 7055
rect -1750 6955 -1745 6995
rect -1705 6955 -1695 6995
rect -1655 6955 -1645 6995
rect -1605 6955 -1595 6995
rect -1555 6955 -1545 6995
rect -1505 6955 -1500 6995
rect -1750 4595 -1500 6955
rect -1750 4555 -1745 4595
rect -1705 4555 -1695 4595
rect -1655 4555 -1645 4595
rect -1605 4555 -1595 4595
rect -1555 4555 -1545 4595
rect -1505 4555 -1500 4595
rect -1750 4495 -1500 4555
rect -1750 4455 -1745 4495
rect -1705 4455 -1695 4495
rect -1655 4455 -1645 4495
rect -1605 4455 -1595 4495
rect -1555 4455 -1545 4495
rect -1505 4455 -1500 4495
rect -1750 4395 -1500 4455
rect -1750 4355 -1745 4395
rect -1705 4355 -1695 4395
rect -1655 4355 -1645 4395
rect -1605 4355 -1595 4395
rect -1555 4355 -1545 4395
rect -1505 4355 -1500 4395
rect -1750 4295 -1500 4355
rect -1750 4255 -1745 4295
rect -1705 4255 -1695 4295
rect -1655 4255 -1645 4295
rect -1605 4255 -1595 4295
rect -1555 4255 -1545 4295
rect -1505 4255 -1500 4295
rect -1750 4195 -1500 4255
rect -1750 4155 -1745 4195
rect -1705 4155 -1695 4195
rect -1655 4155 -1645 4195
rect -1605 4155 -1595 4195
rect -1555 4155 -1545 4195
rect -1505 4155 -1500 4195
rect -1750 4095 -1500 4155
rect -1750 4055 -1745 4095
rect -1705 4055 -1695 4095
rect -1655 4055 -1645 4095
rect -1605 4055 -1595 4095
rect -1555 4055 -1545 4095
rect -1505 4055 -1500 4095
rect -1750 3995 -1500 4055
rect -1750 3955 -1745 3995
rect -1705 3955 -1695 3995
rect -1655 3955 -1645 3995
rect -1605 3955 -1595 3995
rect -1555 3955 -1545 3995
rect -1505 3955 -1500 3995
rect -1750 3745 -1500 3955
rect -1750 3705 -1745 3745
rect -1705 3705 -1695 3745
rect -1655 3705 -1645 3745
rect -1605 3705 -1595 3745
rect -1555 3705 -1545 3745
rect -1505 3705 -1500 3745
rect -1750 3645 -1500 3705
rect -1750 3605 -1745 3645
rect -1705 3605 -1695 3645
rect -1655 3605 -1645 3645
rect -1605 3605 -1595 3645
rect -1555 3605 -1545 3645
rect -1505 3605 -1500 3645
rect -1750 3545 -1500 3605
rect -1750 3505 -1745 3545
rect -1705 3505 -1695 3545
rect -1655 3505 -1645 3545
rect -1605 3505 -1595 3545
rect -1555 3505 -1545 3545
rect -1505 3505 -1500 3545
rect -1750 3445 -1500 3505
rect -1750 3405 -1745 3445
rect -1705 3405 -1695 3445
rect -1655 3405 -1645 3445
rect -1605 3405 -1595 3445
rect -1555 3405 -1545 3445
rect -1505 3405 -1500 3445
rect -1750 3345 -1500 3405
rect -1750 3305 -1745 3345
rect -1705 3305 -1695 3345
rect -1655 3305 -1645 3345
rect -1605 3305 -1595 3345
rect -1555 3305 -1545 3345
rect -1505 3305 -1500 3345
rect -1750 3245 -1500 3305
rect -1750 3205 -1745 3245
rect -1705 3205 -1695 3245
rect -1655 3205 -1645 3245
rect -1605 3205 -1595 3245
rect -1555 3205 -1545 3245
rect -1505 3205 -1500 3245
rect -1750 3145 -1500 3205
rect -1750 3105 -1745 3145
rect -1705 3105 -1695 3145
rect -1655 3105 -1645 3145
rect -1605 3105 -1595 3145
rect -1555 3105 -1545 3145
rect -1505 3105 -1500 3145
rect -1750 745 -1500 3105
rect -1750 705 -1745 745
rect -1705 705 -1695 745
rect -1655 705 -1645 745
rect -1605 705 -1595 745
rect -1555 705 -1545 745
rect -1505 705 -1500 745
rect -1750 645 -1500 705
rect -1750 605 -1745 645
rect -1705 605 -1695 645
rect -1655 605 -1645 645
rect -1605 605 -1595 645
rect -1555 605 -1545 645
rect -1505 605 -1500 645
rect -1750 545 -1500 605
rect -1750 505 -1745 545
rect -1705 505 -1695 545
rect -1655 505 -1645 545
rect -1605 505 -1595 545
rect -1555 505 -1545 545
rect -1505 505 -1500 545
rect -1750 445 -1500 505
rect -1750 405 -1745 445
rect -1705 405 -1695 445
rect -1655 405 -1645 445
rect -1605 405 -1595 445
rect -1555 405 -1545 445
rect -1505 405 -1500 445
rect -1750 345 -1500 405
rect -1750 305 -1745 345
rect -1705 305 -1695 345
rect -1655 305 -1645 345
rect -1605 305 -1595 345
rect -1555 305 -1545 345
rect -1505 305 -1500 345
rect -1750 245 -1500 305
rect -1750 205 -1745 245
rect -1705 205 -1695 245
rect -1655 205 -1645 245
rect -1605 205 -1595 245
rect -1555 205 -1545 245
rect -1505 205 -1500 245
rect -1750 145 -1500 205
rect -1750 105 -1745 145
rect -1705 105 -1695 145
rect -1655 105 -1645 145
rect -1605 105 -1595 145
rect -1555 105 -1545 145
rect -1505 105 -1500 145
rect -1750 0 -1500 105
rect -1450 6695 -1400 7700
rect -1450 6655 -1445 6695
rect -1405 6655 -1400 6695
rect -1450 6295 -1400 6655
rect -1450 6255 -1445 6295
rect -1405 6255 -1400 6295
rect -1450 6095 -1400 6255
rect -1450 6055 -1445 6095
rect -1405 6055 -1400 6095
rect -1450 5895 -1400 6055
rect -1450 5855 -1445 5895
rect -1405 5855 -1400 5895
rect -1450 5695 -1400 5855
rect -1450 5655 -1445 5695
rect -1405 5655 -1400 5695
rect -1450 5495 -1400 5655
rect -1450 5455 -1445 5495
rect -1405 5455 -1400 5495
rect -1450 5295 -1400 5455
rect -1450 5255 -1445 5295
rect -1405 5255 -1400 5295
rect -1450 4895 -1400 5255
rect -1450 4855 -1445 4895
rect -1405 4855 -1400 4895
rect -1450 2845 -1400 4855
rect -1450 2805 -1445 2845
rect -1405 2805 -1400 2845
rect -1450 2445 -1400 2805
rect -1450 2405 -1445 2445
rect -1405 2405 -1400 2445
rect -1450 2245 -1400 2405
rect -1450 2205 -1445 2245
rect -1405 2205 -1400 2245
rect -1450 2045 -1400 2205
rect -1450 2005 -1445 2045
rect -1405 2005 -1400 2045
rect -1450 1845 -1400 2005
rect -1450 1805 -1445 1845
rect -1405 1805 -1400 1845
rect -1450 1645 -1400 1805
rect -1450 1605 -1445 1645
rect -1405 1605 -1400 1645
rect -1450 1445 -1400 1605
rect -1450 1405 -1445 1445
rect -1405 1405 -1400 1445
rect -1450 1045 -1400 1405
rect -1450 1005 -1445 1045
rect -1405 1005 -1400 1045
rect -1450 0 -1400 1005
rect -1350 5995 -1300 7700
rect -1350 5955 -1345 5995
rect -1305 5955 -1300 5995
rect -1350 1745 -1300 5955
rect -1350 1705 -1345 1745
rect -1305 1705 -1300 1745
rect -1350 0 -1300 1705
rect -1250 6695 -1200 7700
rect -1250 6655 -1245 6695
rect -1205 6655 -1200 6695
rect -1250 6295 -1200 6655
rect -1250 6255 -1245 6295
rect -1205 6255 -1200 6295
rect -1250 6095 -1200 6255
rect -1250 6055 -1245 6095
rect -1205 6055 -1200 6095
rect -1250 5895 -1200 6055
rect -1250 5855 -1245 5895
rect -1205 5855 -1200 5895
rect -1250 5695 -1200 5855
rect -1250 5655 -1245 5695
rect -1205 5655 -1200 5695
rect -1250 5495 -1200 5655
rect -1250 5455 -1245 5495
rect -1205 5455 -1200 5495
rect -1250 5295 -1200 5455
rect -1250 5255 -1245 5295
rect -1205 5255 -1200 5295
rect -1250 4895 -1200 5255
rect -1250 4855 -1245 4895
rect -1205 4855 -1200 4895
rect -1250 2845 -1200 4855
rect -1250 2805 -1245 2845
rect -1205 2805 -1200 2845
rect -1250 2445 -1200 2805
rect -1250 2405 -1245 2445
rect -1205 2405 -1200 2445
rect -1250 2245 -1200 2405
rect -1250 2205 -1245 2245
rect -1205 2205 -1200 2245
rect -1250 2045 -1200 2205
rect -1250 2005 -1245 2045
rect -1205 2005 -1200 2045
rect -1250 1845 -1200 2005
rect -1250 1805 -1245 1845
rect -1205 1805 -1200 1845
rect -1250 1645 -1200 1805
rect -1250 1605 -1245 1645
rect -1205 1605 -1200 1645
rect -1250 1445 -1200 1605
rect -1250 1405 -1245 1445
rect -1205 1405 -1200 1445
rect -1250 1045 -1200 1405
rect -1250 1005 -1245 1045
rect -1205 1005 -1200 1045
rect -1250 0 -1200 1005
rect -1150 5595 -1100 7700
rect -1150 5555 -1145 5595
rect -1105 5555 -1100 5595
rect -1150 2145 -1100 5555
rect -1150 2105 -1145 2145
rect -1105 2105 -1100 2145
rect -1150 0 -1100 2105
rect -1050 6695 -1000 7700
rect -1050 6655 -1045 6695
rect -1005 6655 -1000 6695
rect -1050 6295 -1000 6655
rect -1050 6255 -1045 6295
rect -1005 6255 -1000 6295
rect -1050 6095 -1000 6255
rect -1050 6055 -1045 6095
rect -1005 6055 -1000 6095
rect -1050 5895 -1000 6055
rect -1050 5855 -1045 5895
rect -1005 5855 -1000 5895
rect -1050 5695 -1000 5855
rect -1050 5655 -1045 5695
rect -1005 5655 -1000 5695
rect -1050 5495 -1000 5655
rect -1050 5455 -1045 5495
rect -1005 5455 -1000 5495
rect -1050 5295 -1000 5455
rect -1050 5255 -1045 5295
rect -1005 5255 -1000 5295
rect -1050 4895 -1000 5255
rect -1050 4855 -1045 4895
rect -1005 4855 -1000 4895
rect -1050 2845 -1000 4855
rect -1050 2805 -1045 2845
rect -1005 2805 -1000 2845
rect -1050 2445 -1000 2805
rect -1050 2405 -1045 2445
rect -1005 2405 -1000 2445
rect -1050 2245 -1000 2405
rect -1050 2205 -1045 2245
rect -1005 2205 -1000 2245
rect -1050 2045 -1000 2205
rect -1050 2005 -1045 2045
rect -1005 2005 -1000 2045
rect -1050 1845 -1000 2005
rect -1050 1805 -1045 1845
rect -1005 1805 -1000 1845
rect -1050 1645 -1000 1805
rect -1050 1605 -1045 1645
rect -1005 1605 -1000 1645
rect -1050 1445 -1000 1605
rect -1050 1405 -1045 1445
rect -1005 1405 -1000 1445
rect -1050 1045 -1000 1405
rect -1050 1005 -1045 1045
rect -1005 1005 -1000 1045
rect -1050 0 -1000 1005
rect -950 6195 -900 7700
rect -950 6155 -945 6195
rect -905 6155 -900 6195
rect -950 1545 -900 6155
rect -950 1505 -945 1545
rect -905 1505 -900 1545
rect -950 0 -900 1505
rect -850 6695 -800 7700
rect -850 6655 -845 6695
rect -805 6655 -800 6695
rect -850 6295 -800 6655
rect -850 6255 -845 6295
rect -805 6255 -800 6295
rect -850 6095 -800 6255
rect -850 6055 -845 6095
rect -805 6055 -800 6095
rect -850 5895 -800 6055
rect -850 5855 -845 5895
rect -805 5855 -800 5895
rect -850 5695 -800 5855
rect -850 5655 -845 5695
rect -805 5655 -800 5695
rect -850 5495 -800 5655
rect -850 5455 -845 5495
rect -805 5455 -800 5495
rect -850 5295 -800 5455
rect -850 5255 -845 5295
rect -805 5255 -800 5295
rect -850 4895 -800 5255
rect -850 4855 -845 4895
rect -805 4855 -800 4895
rect -850 2845 -800 4855
rect -850 2805 -845 2845
rect -805 2805 -800 2845
rect -850 2445 -800 2805
rect -850 2405 -845 2445
rect -805 2405 -800 2445
rect -850 2245 -800 2405
rect -850 2205 -845 2245
rect -805 2205 -800 2245
rect -850 2045 -800 2205
rect -850 2005 -845 2045
rect -805 2005 -800 2045
rect -850 1845 -800 2005
rect -850 1805 -845 1845
rect -805 1805 -800 1845
rect -850 1645 -800 1805
rect -850 1605 -845 1645
rect -805 1605 -800 1645
rect -850 1445 -800 1605
rect -850 1405 -845 1445
rect -805 1405 -800 1445
rect -850 1045 -800 1405
rect -850 1005 -845 1045
rect -805 1005 -800 1045
rect -850 0 -800 1005
rect -750 5395 -700 7700
rect -750 5355 -745 5395
rect -705 5355 -700 5395
rect -750 2345 -700 5355
rect -750 2305 -745 2345
rect -705 2305 -700 2345
rect -750 0 -700 2305
rect -650 6695 -600 7700
rect -650 6655 -645 6695
rect -605 6655 -600 6695
rect -650 6295 -600 6655
rect -650 6255 -645 6295
rect -605 6255 -600 6295
rect -650 6095 -600 6255
rect -650 6055 -645 6095
rect -605 6055 -600 6095
rect -650 5895 -600 6055
rect -650 5855 -645 5895
rect -605 5855 -600 5895
rect -650 5695 -600 5855
rect -650 5655 -645 5695
rect -605 5655 -600 5695
rect -650 5495 -600 5655
rect -650 5455 -645 5495
rect -605 5455 -600 5495
rect -650 5295 -600 5455
rect -650 5255 -645 5295
rect -605 5255 -600 5295
rect -650 4895 -600 5255
rect -650 4855 -645 4895
rect -605 4855 -600 4895
rect -650 2845 -600 4855
rect -650 2805 -645 2845
rect -605 2805 -600 2845
rect -650 2445 -600 2805
rect -650 2405 -645 2445
rect -605 2405 -600 2445
rect -650 2245 -600 2405
rect -650 2205 -645 2245
rect -605 2205 -600 2245
rect -650 2045 -600 2205
rect -650 2005 -645 2045
rect -605 2005 -600 2045
rect -650 1845 -600 2005
rect -650 1805 -645 1845
rect -605 1805 -600 1845
rect -650 1645 -600 1805
rect -650 1605 -645 1645
rect -605 1605 -600 1645
rect -650 1445 -600 1605
rect -650 1405 -645 1445
rect -605 1405 -600 1445
rect -650 1045 -600 1405
rect -650 1005 -645 1045
rect -605 1005 -600 1045
rect -650 0 -600 1005
rect -400 5795 -350 7700
rect -400 5755 -395 5795
rect -355 5755 -350 5795
rect -400 1945 -350 5755
rect -400 1905 -395 1945
rect -355 1905 -350 1945
rect -400 0 -350 1905
rect -250 5795 -200 7700
rect -250 5755 -245 5795
rect -205 5755 -200 5795
rect -250 1945 -200 5755
rect -250 1905 -245 1945
rect -205 1905 -200 1945
rect -250 0 -200 1905
rect 10350 6695 10400 7700
rect 10350 6655 10355 6695
rect 10395 6655 10400 6695
rect 10350 6295 10400 6655
rect 10350 6255 10355 6295
rect 10395 6255 10400 6295
rect 10350 5295 10400 6255
rect 10350 5255 10355 5295
rect 10395 5255 10400 5295
rect 10350 4895 10400 5255
rect 10350 4855 10355 4895
rect 10395 4855 10400 4895
rect 10350 2845 10400 4855
rect 10350 2805 10355 2845
rect 10395 2805 10400 2845
rect 10350 2445 10400 2805
rect 10350 2405 10355 2445
rect 10395 2405 10400 2445
rect 10350 1445 10400 2405
rect 10350 1405 10355 1445
rect 10395 1405 10400 1445
rect 10350 1045 10400 1405
rect 10350 1005 10355 1045
rect 10395 1005 10400 1045
rect 10350 0 10400 1005
rect 10450 6595 10500 7700
rect 10450 6555 10455 6595
rect 10495 6555 10500 6595
rect 10450 6395 10500 6555
rect 10450 6355 10455 6395
rect 10495 6355 10500 6395
rect 10450 1345 10500 6355
rect 10450 1305 10455 1345
rect 10495 1305 10500 1345
rect 10450 1145 10500 1305
rect 10450 1105 10455 1145
rect 10495 1105 10500 1145
rect 10450 0 10500 1105
rect 10550 6495 10600 7700
rect 10550 6455 10555 6495
rect 10595 6455 10600 6495
rect 10550 1245 10600 6455
rect 10550 1205 10555 1245
rect 10595 1205 10600 1245
rect 10550 0 10600 1205
rect 10650 6595 10700 7700
rect 10650 6555 10655 6595
rect 10695 6555 10700 6595
rect 10650 6395 10700 6555
rect 10650 6355 10655 6395
rect 10695 6355 10700 6395
rect 10650 1345 10700 6355
rect 10650 1305 10655 1345
rect 10695 1305 10700 1345
rect 10650 1145 10700 1305
rect 10650 1105 10655 1145
rect 10695 1105 10700 1145
rect 10650 0 10700 1105
rect 10750 6695 10800 7700
rect 10750 6655 10755 6695
rect 10795 6655 10800 6695
rect 10750 6295 10800 6655
rect 10750 6255 10755 6295
rect 10795 6255 10800 6295
rect 10750 5295 10800 6255
rect 10750 5255 10755 5295
rect 10795 5255 10800 5295
rect 10750 4895 10800 5255
rect 10750 4855 10755 4895
rect 10795 4855 10800 4895
rect 10750 2845 10800 4855
rect 10750 2805 10755 2845
rect 10795 2805 10800 2845
rect 10750 2445 10800 2805
rect 10750 2405 10755 2445
rect 10795 2405 10800 2445
rect 10750 1445 10800 2405
rect 10750 1405 10755 1445
rect 10795 1405 10800 1445
rect 10750 1045 10800 1405
rect 10750 1005 10755 1045
rect 10795 1005 10800 1045
rect 10750 0 10800 1005
rect 10850 5195 10900 7700
rect 10850 5155 10855 5195
rect 10895 5155 10900 5195
rect 10850 4995 10900 5155
rect 10850 4955 10855 4995
rect 10895 4955 10900 4995
rect 10850 2745 10900 4955
rect 10850 2705 10855 2745
rect 10895 2705 10900 2745
rect 10850 2545 10900 2705
rect 10850 2505 10855 2545
rect 10895 2505 10900 2545
rect 10850 0 10900 2505
rect 10950 5095 11000 7700
rect 10950 5055 10955 5095
rect 10995 5055 11000 5095
rect 10950 2645 11000 5055
rect 10950 2605 10955 2645
rect 10995 2605 11000 2645
rect 10950 0 11000 2605
rect 11050 5195 11100 7700
rect 11050 5155 11055 5195
rect 11095 5155 11100 5195
rect 11050 4995 11100 5155
rect 11050 4955 11055 4995
rect 11095 4955 11100 4995
rect 11050 2745 11100 4955
rect 11050 2705 11055 2745
rect 11095 2705 11100 2745
rect 11050 2545 11100 2705
rect 11050 2505 11055 2545
rect 11095 2505 11100 2545
rect 11050 0 11100 2505
rect 11150 6695 11200 7700
rect 11150 6655 11155 6695
rect 11195 6655 11200 6695
rect 11150 6295 11200 6655
rect 11150 6255 11155 6295
rect 11195 6255 11200 6295
rect 11150 5295 11200 6255
rect 11150 5255 11155 5295
rect 11195 5255 11200 5295
rect 11150 4895 11200 5255
rect 11150 4855 11155 4895
rect 11195 4855 11200 4895
rect 11150 2845 11200 4855
rect 11150 2805 11155 2845
rect 11195 2805 11200 2845
rect 11150 2445 11200 2805
rect 11150 2405 11155 2445
rect 11195 2405 11200 2445
rect 11150 1445 11200 2405
rect 11150 1405 11155 1445
rect 11195 1405 11200 1445
rect 11150 1045 11200 1405
rect 11150 1005 11155 1045
rect 11195 1005 11200 1045
rect 11150 0 11200 1005
rect 11250 7595 11500 7700
rect 11250 7555 11255 7595
rect 11295 7555 11305 7595
rect 11345 7555 11355 7595
rect 11395 7555 11405 7595
rect 11445 7555 11455 7595
rect 11495 7555 11500 7595
rect 11250 7495 11500 7555
rect 11250 7455 11255 7495
rect 11295 7455 11305 7495
rect 11345 7455 11355 7495
rect 11395 7455 11405 7495
rect 11445 7455 11455 7495
rect 11495 7455 11500 7495
rect 11250 7395 11500 7455
rect 11250 7355 11255 7395
rect 11295 7355 11305 7395
rect 11345 7355 11355 7395
rect 11395 7355 11405 7395
rect 11445 7355 11455 7395
rect 11495 7355 11500 7395
rect 11250 7295 11500 7355
rect 11250 7255 11255 7295
rect 11295 7255 11305 7295
rect 11345 7255 11355 7295
rect 11395 7255 11405 7295
rect 11445 7255 11455 7295
rect 11495 7255 11500 7295
rect 11250 7195 11500 7255
rect 11250 7155 11255 7195
rect 11295 7155 11305 7195
rect 11345 7155 11355 7195
rect 11395 7155 11405 7195
rect 11445 7155 11455 7195
rect 11495 7155 11500 7195
rect 11250 7095 11500 7155
rect 11250 7055 11255 7095
rect 11295 7055 11305 7095
rect 11345 7055 11355 7095
rect 11395 7055 11405 7095
rect 11445 7055 11455 7095
rect 11495 7055 11500 7095
rect 11250 6995 11500 7055
rect 11250 6955 11255 6995
rect 11295 6955 11305 6995
rect 11345 6955 11355 6995
rect 11395 6955 11405 6995
rect 11445 6955 11455 6995
rect 11495 6955 11500 6995
rect 11250 4595 11500 6955
rect 11250 4555 11255 4595
rect 11295 4555 11305 4595
rect 11345 4555 11355 4595
rect 11395 4555 11405 4595
rect 11445 4555 11455 4595
rect 11495 4555 11500 4595
rect 11250 4495 11500 4555
rect 11250 4455 11255 4495
rect 11295 4455 11305 4495
rect 11345 4455 11355 4495
rect 11395 4455 11405 4495
rect 11445 4455 11455 4495
rect 11495 4455 11500 4495
rect 11250 4395 11500 4455
rect 11250 4355 11255 4395
rect 11295 4355 11305 4395
rect 11345 4355 11355 4395
rect 11395 4355 11405 4395
rect 11445 4355 11455 4395
rect 11495 4355 11500 4395
rect 11250 4295 11500 4355
rect 11250 4255 11255 4295
rect 11295 4255 11305 4295
rect 11345 4255 11355 4295
rect 11395 4255 11405 4295
rect 11445 4255 11455 4295
rect 11495 4255 11500 4295
rect 11250 4195 11500 4255
rect 11250 4155 11255 4195
rect 11295 4155 11305 4195
rect 11345 4155 11355 4195
rect 11395 4155 11405 4195
rect 11445 4155 11455 4195
rect 11495 4155 11500 4195
rect 11250 4095 11500 4155
rect 11250 4055 11255 4095
rect 11295 4055 11305 4095
rect 11345 4055 11355 4095
rect 11395 4055 11405 4095
rect 11445 4055 11455 4095
rect 11495 4055 11500 4095
rect 11250 3995 11500 4055
rect 11250 3955 11255 3995
rect 11295 3955 11305 3995
rect 11345 3955 11355 3995
rect 11395 3955 11405 3995
rect 11445 3955 11455 3995
rect 11495 3955 11500 3995
rect 11250 3745 11500 3955
rect 11250 3705 11255 3745
rect 11295 3705 11305 3745
rect 11345 3705 11355 3745
rect 11395 3705 11405 3745
rect 11445 3705 11455 3745
rect 11495 3705 11500 3745
rect 11250 3645 11500 3705
rect 11250 3605 11255 3645
rect 11295 3605 11305 3645
rect 11345 3605 11355 3645
rect 11395 3605 11405 3645
rect 11445 3605 11455 3645
rect 11495 3605 11500 3645
rect 11250 3545 11500 3605
rect 11250 3505 11255 3545
rect 11295 3505 11305 3545
rect 11345 3505 11355 3545
rect 11395 3505 11405 3545
rect 11445 3505 11455 3545
rect 11495 3505 11500 3545
rect 11250 3445 11500 3505
rect 11250 3405 11255 3445
rect 11295 3405 11305 3445
rect 11345 3405 11355 3445
rect 11395 3405 11405 3445
rect 11445 3405 11455 3445
rect 11495 3405 11500 3445
rect 11250 3345 11500 3405
rect 11250 3305 11255 3345
rect 11295 3305 11305 3345
rect 11345 3305 11355 3345
rect 11395 3305 11405 3345
rect 11445 3305 11455 3345
rect 11495 3305 11500 3345
rect 11250 3245 11500 3305
rect 11250 3205 11255 3245
rect 11295 3205 11305 3245
rect 11345 3205 11355 3245
rect 11395 3205 11405 3245
rect 11445 3205 11455 3245
rect 11495 3205 11500 3245
rect 11250 3145 11500 3205
rect 11250 3105 11255 3145
rect 11295 3105 11305 3145
rect 11345 3105 11355 3145
rect 11395 3105 11405 3145
rect 11445 3105 11455 3145
rect 11495 3105 11500 3145
rect 11250 745 11500 3105
rect 11250 705 11255 745
rect 11295 705 11305 745
rect 11345 705 11355 745
rect 11395 705 11405 745
rect 11445 705 11455 745
rect 11495 705 11500 745
rect 11250 645 11500 705
rect 11250 605 11255 645
rect 11295 605 11305 645
rect 11345 605 11355 645
rect 11395 605 11405 645
rect 11445 605 11455 645
rect 11495 605 11500 645
rect 11250 545 11500 605
rect 11250 505 11255 545
rect 11295 505 11305 545
rect 11345 505 11355 545
rect 11395 505 11405 545
rect 11445 505 11455 545
rect 11495 505 11500 545
rect 11250 445 11500 505
rect 11250 405 11255 445
rect 11295 405 11305 445
rect 11345 405 11355 445
rect 11395 405 11405 445
rect 11445 405 11455 445
rect 11495 405 11500 445
rect 11250 345 11500 405
rect 11250 305 11255 345
rect 11295 305 11305 345
rect 11345 305 11355 345
rect 11395 305 11405 345
rect 11445 305 11455 345
rect 11495 305 11500 345
rect 11250 245 11500 305
rect 11250 205 11255 245
rect 11295 205 11305 245
rect 11345 205 11355 245
rect 11395 205 11405 245
rect 11445 205 11455 245
rect 11495 205 11500 245
rect 11250 145 11500 205
rect 11250 105 11255 145
rect 11295 105 11305 145
rect 11345 105 11355 145
rect 11395 105 11405 145
rect 11445 105 11455 145
rect 11495 105 11500 145
rect 11250 0 11500 105
rect 11550 5800 11600 7700
rect 11650 7550 16750 7650
rect 11650 6750 11750 7550
rect 16650 6750 16750 7550
rect 11650 6595 16750 6750
rect 11650 6555 11655 6595
rect 11695 6555 11705 6595
rect 11745 6555 11755 6595
rect 11795 6555 11805 6595
rect 11845 6555 11855 6595
rect 11895 6555 16605 6595
rect 16645 6555 16655 6595
rect 16695 6555 16705 6595
rect 16745 6555 16750 6595
rect 11650 6550 16750 6555
rect 16800 7645 16950 7650
rect 16800 7605 16805 7645
rect 16845 7605 16905 7645
rect 16945 7605 16950 7645
rect 16800 7595 16950 7605
rect 16800 7555 16805 7595
rect 16845 7555 16905 7595
rect 16945 7555 16950 7595
rect 16800 7545 16950 7555
rect 16800 7505 16805 7545
rect 16845 7505 16905 7545
rect 16945 7505 16950 7545
rect 16800 7495 16950 7505
rect 16800 7455 16805 7495
rect 16845 7455 16905 7495
rect 16945 7455 16950 7495
rect 16800 7445 16950 7455
rect 16800 7405 16805 7445
rect 16845 7405 16905 7445
rect 16945 7405 16950 7445
rect 16800 7395 16950 7405
rect 16800 7355 16805 7395
rect 16845 7355 16905 7395
rect 16945 7355 16950 7395
rect 16800 7345 16950 7355
rect 16800 7305 16805 7345
rect 16845 7305 16905 7345
rect 16945 7305 16950 7345
rect 16800 7295 16950 7305
rect 16800 7255 16805 7295
rect 16845 7255 16905 7295
rect 16945 7255 16950 7295
rect 16800 7245 16950 7255
rect 16800 7205 16805 7245
rect 16845 7205 16905 7245
rect 16945 7205 16950 7245
rect 16800 7195 16950 7205
rect 16800 7155 16805 7195
rect 16845 7155 16905 7195
rect 16945 7155 16950 7195
rect 16800 7145 16950 7155
rect 16800 7105 16805 7145
rect 16845 7105 16905 7145
rect 16945 7105 16950 7145
rect 16800 7095 16950 7105
rect 16800 7055 16805 7095
rect 16845 7055 16905 7095
rect 16945 7055 16950 7095
rect 16800 7045 16950 7055
rect 16800 7005 16805 7045
rect 16845 7005 16905 7045
rect 16945 7005 16950 7045
rect 16800 6995 16950 7005
rect 16800 6955 16805 6995
rect 16845 6955 16905 6995
rect 16945 6955 16950 6995
rect 16800 6945 16950 6955
rect 16800 6905 16805 6945
rect 16845 6905 16905 6945
rect 16945 6905 16950 6945
rect 16800 6895 16950 6905
rect 16800 6855 16805 6895
rect 16845 6855 16905 6895
rect 16945 6855 16950 6895
rect 16800 6845 16950 6855
rect 16800 6805 16805 6845
rect 16845 6805 16905 6845
rect 16945 6805 16950 6845
rect 16800 6795 16950 6805
rect 16800 6755 16805 6795
rect 16845 6755 16905 6795
rect 16945 6755 16950 6795
rect 16800 6745 16950 6755
rect 16800 6705 16805 6745
rect 16845 6705 16905 6745
rect 16945 6705 16950 6745
rect 16800 6695 16950 6705
rect 16800 6655 16805 6695
rect 16845 6655 16905 6695
rect 16945 6655 16950 6695
rect 16800 6645 16950 6655
rect 16800 6605 16805 6645
rect 16845 6605 16905 6645
rect 16945 6605 16950 6645
rect 16800 6595 16950 6605
rect 16800 6555 16805 6595
rect 16845 6555 16905 6595
rect 16945 6555 16950 6595
rect 16800 6550 16950 6555
rect 16900 6545 16950 6550
rect 16900 6505 16905 6545
rect 16945 6505 16950 6545
rect 16900 6495 16950 6505
rect 16900 6455 16905 6495
rect 16945 6455 16950 6495
rect 16900 6445 16950 6455
rect 16900 6405 16905 6445
rect 16945 6405 16950 6445
rect 16900 6400 16950 6405
rect 11650 6395 16750 6400
rect 11650 6355 11655 6395
rect 11695 6355 11705 6395
rect 11745 6355 11755 6395
rect 11795 6355 11805 6395
rect 11845 6355 11855 6395
rect 11895 6355 16605 6395
rect 16645 6355 16655 6395
rect 16695 6355 16705 6395
rect 16745 6355 16750 6395
rect 11650 6200 16750 6355
rect 11650 5950 11750 6200
rect 16650 5950 16750 6200
rect 11650 5850 16750 5950
rect 16800 6395 16950 6400
rect 16800 6355 16805 6395
rect 16845 6355 16905 6395
rect 16945 6355 16950 6395
rect 16800 6345 16950 6355
rect 16800 6305 16805 6345
rect 16845 6305 16905 6345
rect 16945 6305 16950 6345
rect 16800 6295 16950 6305
rect 16800 6255 16805 6295
rect 16845 6255 16905 6295
rect 16945 6255 16950 6295
rect 16800 6245 16950 6255
rect 16800 6205 16805 6245
rect 16845 6205 16905 6245
rect 16945 6205 16950 6245
rect 16800 6195 16950 6205
rect 16800 6155 16805 6195
rect 16845 6155 16905 6195
rect 16945 6155 16950 6195
rect 16800 6145 16950 6155
rect 16800 6105 16805 6145
rect 16845 6105 16905 6145
rect 16945 6105 16950 6145
rect 16800 6095 16950 6105
rect 16800 6055 16805 6095
rect 16845 6055 16905 6095
rect 16945 6055 16950 6095
rect 16800 6045 16950 6055
rect 16800 6005 16805 6045
rect 16845 6005 16905 6045
rect 16945 6005 16950 6045
rect 16800 5945 16950 6005
rect 16800 5905 16805 5945
rect 16845 5905 16905 5945
rect 16945 5905 16950 5945
rect 16800 5895 16950 5905
rect 16800 5855 16805 5895
rect 16845 5855 16905 5895
rect 16945 5855 16950 5895
rect 16800 5850 16950 5855
rect 11550 5750 16950 5800
rect 11550 3895 11600 5750
rect 11650 5600 16750 5700
rect 11650 5350 11750 5600
rect 16650 5350 16750 5600
rect 11650 5195 16750 5350
rect 11650 5155 11655 5195
rect 11695 5155 11705 5195
rect 11745 5155 11755 5195
rect 11795 5155 11805 5195
rect 11845 5155 11855 5195
rect 11895 5155 16605 5195
rect 16645 5155 16655 5195
rect 16695 5155 16705 5195
rect 16745 5155 16750 5195
rect 11650 5150 16750 5155
rect 16800 5695 16950 5700
rect 16800 5655 16805 5695
rect 16845 5655 16905 5695
rect 16945 5655 16950 5695
rect 16800 5645 16950 5655
rect 16800 5605 16805 5645
rect 16845 5605 16905 5645
rect 16945 5605 16950 5645
rect 16800 5545 16950 5605
rect 16800 5505 16805 5545
rect 16845 5505 16905 5545
rect 16945 5505 16950 5545
rect 16800 5495 16950 5505
rect 16800 5455 16805 5495
rect 16845 5455 16905 5495
rect 16945 5455 16950 5495
rect 16800 5445 16950 5455
rect 16800 5405 16805 5445
rect 16845 5405 16905 5445
rect 16945 5405 16950 5445
rect 16800 5395 16950 5405
rect 16800 5355 16805 5395
rect 16845 5355 16905 5395
rect 16945 5355 16950 5395
rect 16800 5345 16950 5355
rect 16800 5305 16805 5345
rect 16845 5305 16905 5345
rect 16945 5305 16950 5345
rect 16800 5295 16950 5305
rect 16800 5255 16805 5295
rect 16845 5255 16905 5295
rect 16945 5255 16950 5295
rect 16800 5245 16950 5255
rect 16800 5205 16805 5245
rect 16845 5205 16905 5245
rect 16945 5205 16950 5245
rect 16800 5195 16950 5205
rect 16800 5155 16805 5195
rect 16845 5155 16905 5195
rect 16945 5155 16950 5195
rect 16800 5150 16950 5155
rect 16900 5145 16950 5150
rect 16900 5105 16905 5145
rect 16945 5105 16950 5145
rect 16900 5095 16950 5105
rect 16900 5055 16905 5095
rect 16945 5055 16950 5095
rect 16900 5045 16950 5055
rect 16900 5005 16905 5045
rect 16945 5005 16950 5045
rect 16900 5000 16950 5005
rect 11650 4995 16750 5000
rect 11650 4955 11655 4995
rect 11695 4955 11705 4995
rect 11745 4955 11755 4995
rect 11795 4955 11805 4995
rect 11845 4955 11855 4995
rect 11895 4955 16605 4995
rect 16645 4955 16655 4995
rect 16695 4955 16705 4995
rect 16745 4955 16750 4995
rect 11650 4800 16750 4955
rect 11650 4000 11750 4800
rect 16650 4000 16750 4800
rect 11650 3900 16750 4000
rect 16800 4995 16950 5000
rect 16800 4955 16805 4995
rect 16845 4955 16905 4995
rect 16945 4955 16950 4995
rect 16800 4945 16950 4955
rect 16800 4905 16805 4945
rect 16845 4905 16905 4945
rect 16945 4905 16950 4945
rect 16800 4895 16950 4905
rect 16800 4855 16805 4895
rect 16845 4855 16905 4895
rect 16945 4855 16950 4895
rect 16800 4845 16950 4855
rect 16800 4805 16805 4845
rect 16845 4805 16905 4845
rect 16945 4805 16950 4845
rect 16800 4795 16950 4805
rect 16800 4755 16805 4795
rect 16845 4755 16905 4795
rect 16945 4755 16950 4795
rect 16800 4745 16950 4755
rect 16800 4705 16805 4745
rect 16845 4705 16905 4745
rect 16945 4705 16950 4745
rect 16800 4695 16950 4705
rect 16800 4655 16805 4695
rect 16845 4655 16905 4695
rect 16945 4655 16950 4695
rect 16800 4645 16950 4655
rect 16800 4605 16805 4645
rect 16845 4605 16905 4645
rect 16945 4605 16950 4645
rect 16800 4595 16950 4605
rect 16800 4555 16805 4595
rect 16845 4555 16905 4595
rect 16945 4555 16950 4595
rect 16800 4545 16950 4555
rect 16800 4505 16805 4545
rect 16845 4505 16905 4545
rect 16945 4505 16950 4545
rect 16800 4495 16950 4505
rect 16800 4455 16805 4495
rect 16845 4455 16905 4495
rect 16945 4455 16950 4495
rect 16800 4445 16950 4455
rect 16800 4405 16805 4445
rect 16845 4405 16905 4445
rect 16945 4405 16950 4445
rect 16800 4395 16950 4405
rect 16800 4355 16805 4395
rect 16845 4355 16905 4395
rect 16945 4355 16950 4395
rect 16800 4345 16950 4355
rect 16800 4305 16805 4345
rect 16845 4305 16905 4345
rect 16945 4305 16950 4345
rect 16800 4295 16950 4305
rect 16800 4255 16805 4295
rect 16845 4255 16905 4295
rect 16945 4255 16950 4295
rect 16800 4245 16950 4255
rect 16800 4205 16805 4245
rect 16845 4205 16905 4245
rect 16945 4205 16950 4245
rect 16800 4195 16950 4205
rect 16800 4155 16805 4195
rect 16845 4155 16905 4195
rect 16945 4155 16950 4195
rect 16800 4145 16950 4155
rect 16800 4105 16805 4145
rect 16845 4105 16905 4145
rect 16945 4105 16950 4145
rect 16800 4095 16950 4105
rect 16800 4055 16805 4095
rect 16845 4055 16905 4095
rect 16945 4055 16950 4095
rect 16800 4045 16950 4055
rect 16800 4005 16805 4045
rect 16845 4005 16905 4045
rect 16945 4005 16950 4045
rect 16800 3995 16950 4005
rect 16800 3955 16805 3995
rect 16845 3955 16905 3995
rect 16945 3955 16950 3995
rect 16800 3945 16950 3955
rect 16800 3905 16805 3945
rect 16845 3905 16905 3945
rect 16945 3905 16950 3945
rect 16800 3900 16950 3905
rect 11550 3855 11555 3895
rect 11595 3855 11600 3895
rect 11550 3845 11600 3855
rect 11550 3805 11555 3845
rect 11595 3805 11600 3845
rect 11550 1950 11600 3805
rect 11650 3700 16750 3800
rect 11650 2900 11750 3700
rect 16650 2900 16750 3700
rect 11650 2745 16750 2900
rect 11650 2705 11655 2745
rect 11695 2705 11705 2745
rect 11745 2705 11755 2745
rect 11795 2705 11805 2745
rect 11845 2705 11855 2745
rect 11895 2705 16605 2745
rect 16645 2705 16655 2745
rect 16695 2705 16705 2745
rect 16745 2705 16750 2745
rect 11650 2700 16750 2705
rect 16800 3795 16950 3800
rect 16800 3755 16805 3795
rect 16845 3755 16905 3795
rect 16945 3755 16950 3795
rect 16800 3745 16950 3755
rect 16800 3705 16805 3745
rect 16845 3705 16905 3745
rect 16945 3705 16950 3745
rect 16800 3695 16950 3705
rect 16800 3655 16805 3695
rect 16845 3655 16905 3695
rect 16945 3655 16950 3695
rect 16800 3645 16950 3655
rect 16800 3605 16805 3645
rect 16845 3605 16905 3645
rect 16945 3605 16950 3645
rect 16800 3595 16950 3605
rect 16800 3555 16805 3595
rect 16845 3555 16905 3595
rect 16945 3555 16950 3595
rect 16800 3545 16950 3555
rect 16800 3505 16805 3545
rect 16845 3505 16905 3545
rect 16945 3505 16950 3545
rect 16800 3495 16950 3505
rect 16800 3455 16805 3495
rect 16845 3455 16905 3495
rect 16945 3455 16950 3495
rect 16800 3445 16950 3455
rect 16800 3405 16805 3445
rect 16845 3405 16905 3445
rect 16945 3405 16950 3445
rect 16800 3395 16950 3405
rect 16800 3355 16805 3395
rect 16845 3355 16905 3395
rect 16945 3355 16950 3395
rect 16800 3345 16950 3355
rect 16800 3305 16805 3345
rect 16845 3305 16905 3345
rect 16945 3305 16950 3345
rect 16800 3295 16950 3305
rect 16800 3255 16805 3295
rect 16845 3255 16905 3295
rect 16945 3255 16950 3295
rect 16800 3245 16950 3255
rect 16800 3205 16805 3245
rect 16845 3205 16905 3245
rect 16945 3205 16950 3245
rect 16800 3195 16950 3205
rect 16800 3155 16805 3195
rect 16845 3155 16905 3195
rect 16945 3155 16950 3195
rect 16800 3145 16950 3155
rect 16800 3105 16805 3145
rect 16845 3105 16905 3145
rect 16945 3105 16950 3145
rect 16800 3095 16950 3105
rect 16800 3055 16805 3095
rect 16845 3055 16905 3095
rect 16945 3055 16950 3095
rect 16800 3045 16950 3055
rect 16800 3005 16805 3045
rect 16845 3005 16905 3045
rect 16945 3005 16950 3045
rect 16800 2995 16950 3005
rect 16800 2955 16805 2995
rect 16845 2955 16905 2995
rect 16945 2955 16950 2995
rect 16800 2945 16950 2955
rect 16800 2905 16805 2945
rect 16845 2905 16905 2945
rect 16945 2905 16950 2945
rect 16800 2895 16950 2905
rect 16800 2855 16805 2895
rect 16845 2855 16905 2895
rect 16945 2855 16950 2895
rect 16800 2845 16950 2855
rect 16800 2805 16805 2845
rect 16845 2805 16905 2845
rect 16945 2805 16950 2845
rect 16800 2795 16950 2805
rect 16800 2755 16805 2795
rect 16845 2755 16905 2795
rect 16945 2755 16950 2795
rect 16800 2745 16950 2755
rect 16800 2705 16805 2745
rect 16845 2705 16905 2745
rect 16945 2705 16950 2745
rect 16800 2700 16950 2705
rect 16900 2695 16950 2700
rect 16900 2655 16905 2695
rect 16945 2655 16950 2695
rect 16900 2645 16950 2655
rect 16900 2605 16905 2645
rect 16945 2605 16950 2645
rect 16900 2595 16950 2605
rect 16900 2555 16905 2595
rect 16945 2555 16950 2595
rect 16900 2550 16950 2555
rect 11650 2545 16750 2550
rect 11650 2505 11655 2545
rect 11695 2505 11705 2545
rect 11745 2505 11755 2545
rect 11795 2505 11805 2545
rect 11845 2505 11855 2545
rect 11895 2505 16605 2545
rect 16645 2505 16655 2545
rect 16695 2505 16705 2545
rect 16745 2505 16750 2545
rect 11650 2350 16750 2505
rect 11650 2100 11750 2350
rect 16650 2100 16750 2350
rect 11650 2000 16750 2100
rect 16800 2545 16950 2550
rect 16800 2505 16805 2545
rect 16845 2505 16905 2545
rect 16945 2505 16950 2545
rect 16800 2495 16950 2505
rect 16800 2455 16805 2495
rect 16845 2455 16905 2495
rect 16945 2455 16950 2495
rect 16800 2445 16950 2455
rect 16800 2405 16805 2445
rect 16845 2405 16905 2445
rect 16945 2405 16950 2445
rect 16800 2395 16950 2405
rect 16800 2355 16805 2395
rect 16845 2355 16905 2395
rect 16945 2355 16950 2395
rect 16800 2345 16950 2355
rect 16800 2305 16805 2345
rect 16845 2305 16905 2345
rect 16945 2305 16950 2345
rect 16800 2295 16950 2305
rect 16800 2255 16805 2295
rect 16845 2255 16905 2295
rect 16945 2255 16950 2295
rect 16800 2245 16950 2255
rect 16800 2205 16805 2245
rect 16845 2205 16905 2245
rect 16945 2205 16950 2245
rect 16800 2195 16950 2205
rect 16800 2155 16805 2195
rect 16845 2155 16905 2195
rect 16945 2155 16950 2195
rect 16800 2145 16950 2155
rect 16800 2105 16805 2145
rect 16845 2105 16905 2145
rect 16945 2105 16950 2145
rect 16800 2095 16950 2105
rect 16800 2055 16805 2095
rect 16845 2055 16905 2095
rect 16945 2055 16950 2095
rect 16800 2045 16950 2055
rect 16800 2005 16805 2045
rect 16845 2005 16905 2045
rect 16945 2005 16950 2045
rect 16800 2000 16950 2005
rect 11550 1900 16950 1950
rect 11550 0 11600 1900
rect 11650 1750 16750 1850
rect 11650 1500 11750 1750
rect 16650 1500 16750 1750
rect 11650 1345 16750 1500
rect 11650 1305 11655 1345
rect 11695 1305 11705 1345
rect 11745 1305 11755 1345
rect 11795 1305 11805 1345
rect 11845 1305 11855 1345
rect 11895 1305 16605 1345
rect 16645 1305 16655 1345
rect 16695 1305 16705 1345
rect 16745 1305 16750 1345
rect 11650 1300 16750 1305
rect 16800 1845 16950 1850
rect 16800 1805 16805 1845
rect 16845 1805 16905 1845
rect 16945 1805 16950 1845
rect 16800 1795 16950 1805
rect 16800 1755 16805 1795
rect 16845 1755 16905 1795
rect 16945 1755 16950 1795
rect 16800 1745 16950 1755
rect 16800 1705 16805 1745
rect 16845 1705 16905 1745
rect 16945 1705 16950 1745
rect 16800 1695 16950 1705
rect 16800 1655 16805 1695
rect 16845 1655 16905 1695
rect 16945 1655 16950 1695
rect 16800 1645 16950 1655
rect 16800 1605 16805 1645
rect 16845 1605 16905 1645
rect 16945 1605 16950 1645
rect 16800 1595 16950 1605
rect 16800 1555 16805 1595
rect 16845 1555 16905 1595
rect 16945 1555 16950 1595
rect 16800 1545 16950 1555
rect 16800 1505 16805 1545
rect 16845 1505 16905 1545
rect 16945 1505 16950 1545
rect 16800 1495 16950 1505
rect 16800 1455 16805 1495
rect 16845 1455 16905 1495
rect 16945 1455 16950 1495
rect 16800 1445 16950 1455
rect 16800 1405 16805 1445
rect 16845 1405 16905 1445
rect 16945 1405 16950 1445
rect 16800 1395 16950 1405
rect 16800 1355 16805 1395
rect 16845 1355 16905 1395
rect 16945 1355 16950 1395
rect 16800 1345 16950 1355
rect 16800 1305 16805 1345
rect 16845 1305 16905 1345
rect 16945 1305 16950 1345
rect 16800 1300 16950 1305
rect 16900 1295 16950 1300
rect 16900 1255 16905 1295
rect 16945 1255 16950 1295
rect 16900 1245 16950 1255
rect 16900 1205 16905 1245
rect 16945 1205 16950 1245
rect 16900 1195 16950 1205
rect 16900 1155 16905 1195
rect 16945 1155 16950 1195
rect 16900 1150 16950 1155
rect 11650 1145 16750 1150
rect 11650 1105 11655 1145
rect 11695 1105 11705 1145
rect 11745 1105 11755 1145
rect 11795 1105 11805 1145
rect 11845 1105 11855 1145
rect 11895 1105 16605 1145
rect 16645 1105 16655 1145
rect 16695 1105 16705 1145
rect 16745 1105 16750 1145
rect 11650 950 16750 1105
rect 11650 150 11750 950
rect 16650 150 16750 950
rect 11650 50 16750 150
rect 16800 1145 16950 1150
rect 16800 1105 16805 1145
rect 16845 1105 16905 1145
rect 16945 1105 16950 1145
rect 16800 1095 16950 1105
rect 16800 1055 16805 1095
rect 16845 1055 16905 1095
rect 16945 1055 16950 1095
rect 16800 1045 16950 1055
rect 16800 1005 16805 1045
rect 16845 1005 16905 1045
rect 16945 1005 16950 1045
rect 16800 995 16950 1005
rect 16800 955 16805 995
rect 16845 955 16905 995
rect 16945 955 16950 995
rect 16800 945 16950 955
rect 16800 905 16805 945
rect 16845 905 16905 945
rect 16945 905 16950 945
rect 16800 895 16950 905
rect 16800 855 16805 895
rect 16845 855 16905 895
rect 16945 855 16950 895
rect 16800 845 16950 855
rect 16800 805 16805 845
rect 16845 805 16905 845
rect 16945 805 16950 845
rect 16800 795 16950 805
rect 16800 755 16805 795
rect 16845 755 16905 795
rect 16945 755 16950 795
rect 16800 745 16950 755
rect 16800 705 16805 745
rect 16845 705 16905 745
rect 16945 705 16950 745
rect 16800 695 16950 705
rect 16800 655 16805 695
rect 16845 655 16905 695
rect 16945 655 16950 695
rect 16800 645 16950 655
rect 16800 605 16805 645
rect 16845 605 16905 645
rect 16945 605 16950 645
rect 16800 595 16950 605
rect 16800 555 16805 595
rect 16845 555 16905 595
rect 16945 555 16950 595
rect 16800 545 16950 555
rect 16800 505 16805 545
rect 16845 505 16905 545
rect 16945 505 16950 545
rect 16800 495 16950 505
rect 16800 455 16805 495
rect 16845 455 16905 495
rect 16945 455 16950 495
rect 16800 445 16950 455
rect 16800 405 16805 445
rect 16845 405 16905 445
rect 16945 405 16950 445
rect 16800 395 16950 405
rect 16800 355 16805 395
rect 16845 355 16905 395
rect 16945 355 16950 395
rect 16800 345 16950 355
rect 16800 305 16805 345
rect 16845 305 16905 345
rect 16945 305 16950 345
rect 16800 295 16950 305
rect 16800 255 16805 295
rect 16845 255 16905 295
rect 16945 255 16950 295
rect 16800 245 16950 255
rect 16800 205 16805 245
rect 16845 205 16905 245
rect 16945 205 16950 245
rect 16800 195 16950 205
rect 16800 155 16805 195
rect 16845 155 16905 195
rect 16945 155 16950 195
rect 16800 145 16950 155
rect 16800 105 16805 145
rect 16845 105 16905 145
rect 16945 105 16950 145
rect 16800 95 16950 105
rect 16800 55 16805 95
rect 16845 55 16905 95
rect 16945 55 16950 95
rect 16800 50 16950 55
use ddac_slice  ddab_slice_0
timestamp 1723498139
transform 1 0 3200 0 1 0
box -3200 0 6550 3850
use ddac_slice  ddab_slice_1
timestamp 1723498139
transform -1 0 6550 0 -1 7700
box -3200 0 6550 3850
use invdummy  invdummy_0
timestamp 1722856725
transform -1 0 9900 0 -1 7700
box -50 0 300 3850
use invdummy  invdummy_1
timestamp 1722856725
transform 1 0 -150 0 -1 7700
box -50 0 300 3850
use invdummy  invdummy_2
timestamp 1722856725
transform -1 0 9900 0 1 0
box -50 0 300 3850
use invdummy  invdummy_3
timestamp 1722856725
transform 1 0 -150 0 1 0
box -50 0 300 3850
use invedge  invedge_0
timestamp 1722865417
transform 1 0 9700 0 -1 8800
box 150 1100 600 4950
use invedge  invedge_1
timestamp 1722865417
transform -1 0 50 0 -1 8800
box 150 1100 600 4950
use invedge  invedge_2
timestamp 1722865417
transform 1 0 9700 0 1 -1100
box 150 1100 600 4950
use invedge  invedge_3
timestamp 1722865417
transform -1 0 50 0 1 -1100
box 150 1100 600 4950
<< labels >>
rlabel metal4 -1350 7650 -1300 7700 0 ipa
port 1 nsew
rlabel metal4 -1150 7650 -1100 7700 0 ima
port 2 nsew
rlabel metal4 -950 7650 -900 7700 0 ipb
port 3 nsew
rlabel metal4 -750 7650 -700 7700 0 imb
port 4 nsew
rlabel metal4 10850 7650 10900 7700 0 op
port 5 nsew
rlabel metal4 11050 7650 11100 7700 0 op
port 5 nsew
rlabel metal4 10450 7650 10500 7700 0 om
port 6 nsew
rlabel metal4 10650 7650 10700 7700 0 om
port 6 nsew
rlabel metal4 -400 7650 -350 7700 0 bp
port 7 nsew
rlabel metal4 -250 7650 -200 7700 0 bn
port 8 nsew
rlabel metal4 -1750 7650 -1500 7700 0 vdd
port 9 nsew
rlabel metal4 -1450 7650 -1400 7700 0 vss
port 10 nsew
rlabel metal4 -1850 7650 -1800 7700 0 vsub
port 11 nsew
rlabel metal4 10550 7650 10600 7700 0 xp
rlabel metal4 10950 7650 11000 7700 0 xm
<< end >>
