* NGSPICE file created from ddab_slice0.ext - technology: sky130A

.subckt inv1p1 in out bp bn vreg vss vsub
X0 vreg in out bp sky130_fd_pr__pfet_01v8_lvt ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=4
X1 out in vreg bp sky130_fd_pr__pfet_01v8_lvt ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=4
X2 out in xt bn sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=4
X3 out in xb bn sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=4
X4 out in vreg bp sky130_fd_pr__pfet_01v8_lvt ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=4
X5 xt in vss bn sky130_fd_pr__nfet_01v8 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=4
X6 vreg in out bp sky130_fd_pr__pfet_01v8_lvt ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=4
X7 xb in vss bn sky130_fd_pr__nfet_01v8 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=4
.ends

.subckt ddab_slice0 ip im xm xp op om bp bn vdd vss vsub
Xa0 ip xm bp bn vdd vss vsub inv1p1
Xa1 xp xm bp bn vdd vss vsub inv1p1
Xa2 xm xm bp bn vdd vss vsub inv1p1
Xa3 ip xm bp bn vdd vss vsub inv1p1
Xa4 im xp bp bn vdd vss vsub inv1p1
Xa6 xm xp bp bn vdd vss vsub inv1p1
Xa5 xp xp bp bn vdd vss vsub inv1p1
Xa7 im xp bp bn vdd vss vsub inv1p1
.ends

