magic
tech sky130A
timestamp 1726447784
<< locali >>
rect 50 3800 7300 3850
rect 50 2900 7300 2950
rect 50 2750 7300 2800
rect 4550 1235 4600 1250
rect 4550 1215 4565 1235
rect 4585 1215 4600 1235
rect 4550 1200 4600 1215
rect 50 1050 7300 1100
rect 50 900 7300 950
rect 50 0 7300 50
<< viali >>
rect 4565 1215 4585 1235
<< metal1 >>
rect 6350 1940 6400 1950
rect 6350 1910 6360 1940
rect 6390 1910 6400 1940
rect 6350 1900 6400 1910
rect 4550 1240 4600 1250
rect 4550 1210 4560 1240
rect 4590 1210 4600 1240
rect 4550 1200 4600 1210
<< via1 >>
rect 2760 2610 2790 2640
rect 960 1910 990 1940
rect 6360 1910 6390 1940
rect 4560 1235 4590 1240
rect 4560 1215 4565 1235
rect 4565 1215 4585 1235
rect 4585 1215 4590 1235
rect 4560 1210 4590 1215
<< metal2 >>
rect 2750 2640 2800 2650
rect 2750 2610 2760 2640
rect 2790 2610 2800 2640
rect 2750 2600 2800 2610
rect 950 1940 6400 1950
rect 950 1910 960 1940
rect 990 1910 6360 1940
rect 6390 1910 6400 1940
rect 950 1900 6400 1910
rect 4550 1240 4600 1250
rect 4550 1210 4560 1240
rect 4590 1210 4600 1240
rect 4550 1200 4600 1210
<< via2 >>
rect 2760 2610 2790 2640
rect 4560 1210 4590 1240
<< metal3 >>
rect 50 3700 7300 3750
rect 50 2800 7300 2850
rect 50 2745 7300 2750
rect 50 2705 505 2745
rect 545 2705 7300 2745
rect 50 2700 7300 2705
rect 50 2640 7300 2650
rect 50 2610 2760 2640
rect 2790 2610 7300 2640
rect 50 2600 7300 2610
rect 50 2545 7300 2550
rect 50 2505 505 2545
rect 545 2505 7300 2545
rect 50 2500 7300 2505
rect 50 2100 7300 2150
rect 50 1700 7300 1750
rect 50 1345 7300 1350
rect 50 1305 6805 1345
rect 6845 1305 7300 1345
rect 50 1300 7300 1305
rect 50 1240 7300 1250
rect 50 1210 4560 1240
rect 4590 1210 7300 1240
rect 50 1200 7300 1210
rect 50 1145 7300 1150
rect 50 1105 6805 1145
rect 6845 1105 7300 1145
rect 50 1100 7300 1105
rect 50 1000 7300 1050
rect 50 100 7300 150
<< via3 >>
rect 505 2705 545 2745
rect 505 2505 545 2545
rect 6805 1305 6845 1345
rect 6805 1105 6845 1145
<< metal4 >>
rect 500 2745 550 2750
rect 500 2705 505 2745
rect 545 2705 550 2745
rect 500 2700 550 2705
rect 500 2545 550 2550
rect 500 2505 505 2545
rect 545 2505 550 2545
rect 500 2500 550 2505
rect 6800 1345 6850 1350
rect 6800 1305 6805 1345
rect 6845 1305 6850 1345
rect 6800 1300 6850 1305
rect 6800 1145 6850 1150
rect 6800 1105 6805 1145
rect 6845 1105 6850 1145
rect 6800 1100 6850 1105
use inv1p1  a0
timestamp 1726000395
transform 1 0 50 0 1 0
box -50 0 1000 3850
use inv1p1  a1
timestamp 1726000395
transform -1 0 1900 0 1 0
box -50 0 1000 3850
use inv1p1  a2
timestamp 1726000395
transform 1 0 1850 0 1 0
box -50 0 1000 3850
use inv1p1  a3
timestamp 1726000395
transform -1 0 3700 0 1 0
box -50 0 1000 3850
use inv1p1  a4
timestamp 1726000395
transform 1 0 3650 0 1 0
box -50 0 1000 3850
use inv1p1  a5
timestamp 1726000395
transform -1 0 5500 0 1 0
box -50 0 1000 3850
use inv1p1  a6
timestamp 1726000395
transform 1 0 5450 0 1 0
box -50 0 1000 3850
use inv1p1  a7
timestamp 1726000395
transform -1 0 7300 0 1 0
box -50 0 1000 3850
<< labels >>
rlabel metal3 50 2100 7300 2150 0 ip
port 1 nsew
rlabel metal3 50 1700 7300 1750 0 im
port 2 nsew
rlabel metal3 50 1200 7300 1250 0 xm
port 3 nsew
rlabel metal3 50 2600 7300 2650 0 xp
port 4 nsew
rlabel metal3 50 2700 7300 2750 0 op
port 5 nsew
rlabel metal3 50 2500 7300 2550 0 op
port 5 nsew
rlabel metal3 50 1300 7300 1350 0 om
port 6 nsew
rlabel metal3 50 1100 7300 1150 0 om
port 6 nsew
rlabel locali 50 2900 7300 2950 0 bp
port 7 nsew
rlabel locali 50 900 7300 950 0 bp
port 7 nsew
rlabel locali 50 2750 7300 2800 0 bn
port 8 nsew
rlabel locali 50 1050 7300 1100 0 bn
port 8 nsew
rlabel metal3 50 3700 7300 3750 0 vdd
port 9 nsew
rlabel metal3 50 100 7300 150 0 vdd
port 9 nsew
rlabel metal3 50 2800 7300 2850 0 vss
port 10 nsew
rlabel metal3 50 1000 7300 1050 0 vss
port 10 nsew
rlabel metal2 3650 1900 3700 1950 0 x
rlabel locali 50 3800 7300 3850 0 vsub
port 11 nsew
rlabel locali 50 0 7300 50 0 vsub
port 11 nsew
<< end >>
