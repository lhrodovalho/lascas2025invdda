magic
tech sky130A
timestamp 1726835717
<< dnwell >>
rect -9500 9600 -9450 9650
rect -9350 9600 -9300 9650
<< nwell >>
rect -9500 9600 -9450 9650
<< pwell >>
rect -9350 9600 -9300 9650
<< psubdiff >>
rect -9350 9635 -9300 9650
rect -9350 9615 -9335 9635
rect -9315 9615 -9300 9635
rect -9350 9600 -9300 9615
<< nsubdiff >>
rect -9500 9635 -9450 9650
rect -9500 9615 -9485 9635
rect -9465 9615 -9450 9635
rect -9500 9600 -9450 9615
<< psubdiffcont >>
rect -9335 9615 -9315 9635
<< nsubdiffcont >>
rect -9485 9615 -9465 9635
<< locali >>
rect -9500 13485 -9450 13500
rect -9500 13465 -9485 13485
rect -9465 13465 -9450 13485
rect -9500 13450 -9450 13465
rect -9350 13485 -9300 13500
rect -9350 13465 -9335 13485
rect -9315 13465 -9300 13485
rect -9350 13450 -9300 13465
rect -9650 11585 -9600 11600
rect -9650 11565 -9635 11585
rect -9615 11565 -9600 11585
rect -9650 11535 -9600 11565
rect -9650 11515 -9635 11535
rect -9615 11515 -9600 11535
rect -9650 11500 -9600 11515
rect -9500 9635 -9450 9650
rect -9500 9615 -9485 9635
rect -9465 9615 -9450 9635
rect -9500 9600 -9450 9615
rect -9350 9635 -9300 9650
rect -9350 9615 -9335 9635
rect -9315 9615 -9300 9635
rect -9350 9600 -9300 9615
<< viali >>
rect -9485 13465 -9465 13485
rect -9335 13465 -9315 13485
rect -9635 11565 -9615 11585
rect -9635 11515 -9615 11535
rect -9485 9615 -9465 9635
rect -9335 9615 -9315 9635
<< metal1 >>
rect -9500 13490 -9450 13500
rect -9500 13460 -9490 13490
rect -9460 13460 -9450 13490
rect -9500 13450 -9450 13460
rect -9350 13490 -9300 13500
rect -9350 13460 -9340 13490
rect -9310 13460 -9300 13490
rect -9350 13450 -9300 13460
rect -9650 11590 -9600 11600
rect -9650 11560 -9640 11590
rect -9610 11560 -9600 11590
rect -9650 11540 -9600 11560
rect -9650 11510 -9640 11540
rect -9610 11510 -9600 11540
rect -9650 11500 -9600 11510
rect -9500 9640 -9450 9650
rect -9500 9610 -9490 9640
rect -9460 9610 -9450 9640
rect -9500 9600 -9450 9610
rect -9350 9640 -9300 9650
rect -9350 9610 -9340 9640
rect -9310 9610 -9300 9640
rect -9350 9600 -9300 9610
<< via1 >>
rect -9490 13485 -9460 13490
rect -9490 13465 -9485 13485
rect -9485 13465 -9465 13485
rect -9465 13465 -9460 13485
rect -9490 13460 -9460 13465
rect -9340 13485 -9310 13490
rect -9340 13465 -9335 13485
rect -9335 13465 -9315 13485
rect -9315 13465 -9310 13485
rect -9340 13460 -9310 13465
rect -9640 11585 -9610 11590
rect -9640 11565 -9635 11585
rect -9635 11565 -9615 11585
rect -9615 11565 -9610 11585
rect -9640 11560 -9610 11565
rect -9640 11535 -9610 11540
rect -9640 11515 -9635 11535
rect -9635 11515 -9615 11535
rect -9615 11515 -9610 11535
rect -9640 11510 -9610 11515
rect -9490 9635 -9460 9640
rect -9490 9615 -9485 9635
rect -9485 9615 -9465 9635
rect -9465 9615 -9460 9635
rect -9490 9610 -9460 9615
rect -9340 9635 -9310 9640
rect -9340 9615 -9335 9635
rect -9335 9615 -9315 9635
rect -9315 9615 -9310 9635
rect -9340 9610 -9310 9615
<< metal2 >>
rect -9500 13490 -9450 13500
rect -9500 13460 -9490 13490
rect -9460 13460 -9450 13490
rect -9500 13450 -9450 13460
rect -9350 13490 -9300 13500
rect -9350 13460 -9340 13490
rect -9310 13460 -9300 13490
rect -9350 13450 -9300 13460
rect -10950 11590 13200 11600
rect -10950 11560 -10940 11590
rect -10910 11560 -9640 11590
rect -9610 11560 13200 11590
rect -10950 11540 13200 11560
rect -10950 11510 -10940 11540
rect -10910 11510 -9640 11540
rect -9610 11510 13200 11540
rect -10950 11500 13200 11510
rect -9500 9640 -9450 9650
rect -9500 9610 -9490 9640
rect -9460 9610 -9450 9640
rect -9500 9600 -9450 9610
rect -9350 9640 -9300 9650
rect -9350 9610 -9340 9640
rect -9310 9610 -9300 9640
rect -9350 9600 -9300 9610
<< via2 >>
rect -9490 13460 -9460 13490
rect -9340 13460 -9310 13490
rect -10940 11560 -10910 11590
rect -9640 11560 -9610 11590
rect -10940 11510 -10910 11540
rect -9640 11510 -9610 11540
rect -9490 9610 -9460 9640
rect -9340 9610 -9310 9640
<< metal3 >>
rect 14050 15395 21950 15400
rect 14050 15355 14055 15395
rect 14095 15355 21905 15395
rect 21945 15355 21950 15395
rect 14050 15350 21950 15355
rect -10850 15295 -9650 15300
rect -10850 15255 -10845 15295
rect -10805 15255 -10795 15295
rect -10755 15255 -10745 15295
rect -10705 15255 -10695 15295
rect -10655 15255 -10645 15295
rect -10605 15255 -9650 15295
rect -10850 15250 -9650 15255
rect -10850 15195 -9650 15200
rect -10850 15155 -10845 15195
rect -10805 15155 -10795 15195
rect -10755 15155 -10745 15195
rect -10705 15155 -10695 15195
rect -10655 15155 -10645 15195
rect -10605 15155 -9650 15195
rect -10850 15150 -9650 15155
rect -10850 15095 -9650 15100
rect -10850 15055 -10845 15095
rect -10805 15055 -10795 15095
rect -10755 15055 -10745 15095
rect -10705 15055 -10695 15095
rect -10655 15055 -10645 15095
rect -10605 15055 -9650 15095
rect -10850 15050 -9650 15055
rect -10850 14995 -9650 15000
rect -10850 14955 -10845 14995
rect -10805 14955 -10795 14995
rect -10755 14955 -10745 14995
rect -10705 14955 -10695 14995
rect -10655 14955 -10645 14995
rect -10605 14955 -9650 14995
rect -10850 14950 -9650 14955
rect -10850 14895 -9650 14900
rect -10850 14855 -10845 14895
rect -10805 14855 -10795 14895
rect -10755 14855 -10745 14895
rect -10705 14855 -10695 14895
rect -10655 14855 -10645 14895
rect -10605 14855 -9650 14895
rect -10850 14850 -9650 14855
rect -10850 14795 -9650 14800
rect -10850 14755 -10845 14795
rect -10805 14755 -10795 14795
rect -10755 14755 -10745 14795
rect -10705 14755 -10695 14795
rect -10655 14755 -10645 14795
rect -10605 14755 -9650 14795
rect -10850 14750 -9650 14755
rect -10850 14695 -9650 14700
rect -10850 14655 -10845 14695
rect -10805 14655 -10795 14695
rect -10755 14655 -10745 14695
rect -10705 14655 -10695 14695
rect -10655 14655 -10645 14695
rect -10605 14655 -9650 14695
rect -10850 14650 -9650 14655
rect -10550 14395 -9650 14400
rect -10550 14355 -10545 14395
rect -10505 14355 -10345 14395
rect -10305 14355 -10145 14395
rect -10105 14355 -9945 14395
rect -9905 14355 -9745 14395
rect -9705 14355 -9650 14395
rect -10550 14350 -9650 14355
rect 13200 14395 14100 14400
rect 13200 14355 13255 14395
rect 13295 14355 13655 14395
rect 13695 14355 14100 14395
rect 13200 14350 14100 14355
rect 12600 14295 13600 14300
rect 12600 14255 13355 14295
rect 13395 14255 13555 14295
rect 13595 14255 13600 14295
rect 12600 14250 13600 14255
rect 12600 14195 13500 14200
rect 12600 14155 13455 14195
rect 13495 14155 13500 14195
rect 12600 14150 13500 14155
rect 12600 14095 13600 14100
rect 12600 14055 13355 14095
rect 13395 14055 13555 14095
rect 13595 14055 13600 14095
rect 12600 14050 13600 14055
rect -10550 13995 -9650 14000
rect -10550 13955 -10545 13995
rect -10505 13955 -10345 13995
rect -10305 13955 -10145 13995
rect -10105 13955 -9945 13995
rect -9905 13955 -9745 13995
rect -9705 13955 -9650 13995
rect -10550 13950 -9650 13955
rect 13200 13995 14100 14000
rect 13200 13955 13255 13995
rect 13295 13955 13655 13995
rect 13695 13955 14100 13995
rect 13200 13950 14100 13955
rect -10550 13895 -9650 13900
rect -10550 13855 -10545 13895
rect -10505 13855 -10345 13895
rect -10305 13855 -10145 13895
rect -10105 13855 -9945 13895
rect -9905 13855 -9745 13895
rect -9705 13855 -9650 13895
rect -10550 13850 -9650 13855
rect 13200 13895 14100 13900
rect 13200 13855 13255 13895
rect 13295 13855 13655 13895
rect 13695 13855 14100 13895
rect 13200 13850 14100 13855
rect -10550 13795 -9650 13800
rect -10550 13755 -10545 13795
rect -10505 13755 -10345 13795
rect -10305 13755 -10145 13795
rect -10105 13755 -9945 13795
rect -9905 13755 -9745 13795
rect -9705 13755 -9650 13795
rect -10550 13750 -9650 13755
rect 13200 13795 14100 13800
rect 13200 13755 13255 13795
rect 13295 13755 13655 13795
rect 13695 13755 14100 13795
rect 13200 13750 14100 13755
rect -10250 13695 -9050 13700
rect -10250 13655 -10245 13695
rect -10205 13655 -9050 13695
rect -10250 13650 -9050 13655
rect 13200 13695 14100 13700
rect 13200 13655 13255 13695
rect 13295 13655 13655 13695
rect 13695 13655 14100 13695
rect 13200 13650 14100 13655
rect -10550 13595 -9650 13600
rect -10550 13555 -10545 13595
rect -10505 13555 -10345 13595
rect -10305 13555 -10145 13595
rect -10105 13555 -9945 13595
rect -9905 13555 -9745 13595
rect -9705 13555 -9650 13595
rect -10550 13550 -9650 13555
rect 13200 13595 14100 13600
rect 13200 13555 13255 13595
rect 13295 13555 13655 13595
rect 13695 13555 14100 13595
rect 13200 13550 14100 13555
rect -9500 13495 -9450 13500
rect -9500 13455 -9495 13495
rect -9455 13455 -9450 13495
rect -9500 13450 -9450 13455
rect -9350 13495 -9300 13500
rect -9350 13455 -9345 13495
rect -9305 13455 -9300 13495
rect -9350 13450 -9300 13455
rect -10550 13395 -9650 13400
rect -10550 13355 -10545 13395
rect -10505 13355 -10345 13395
rect -10305 13355 -10145 13395
rect -10105 13355 -9945 13395
rect -9905 13355 -9745 13395
rect -9705 13355 -9650 13395
rect -10550 13350 -9650 13355
rect 13200 13395 14100 13400
rect 13200 13355 13255 13395
rect 13295 13355 13655 13395
rect 13695 13355 14100 13395
rect 13200 13350 14100 13355
rect -10450 13295 -9050 13300
rect -10450 13255 -10445 13295
rect -10405 13255 -9050 13295
rect -10450 13250 -9050 13255
rect 13200 13295 14100 13300
rect 13200 13255 13255 13295
rect 13295 13255 13655 13295
rect 13695 13255 14100 13295
rect 13200 13250 14100 13255
rect -10550 13195 -9650 13200
rect -10550 13155 -10545 13195
rect -10505 13155 -10345 13195
rect -10305 13155 -10145 13195
rect -10105 13155 -9945 13195
rect -9905 13155 -9745 13195
rect -9705 13155 -9650 13195
rect -10550 13150 -9650 13155
rect 13200 13195 14100 13200
rect 13200 13155 13255 13195
rect 13295 13155 13655 13195
rect 13695 13155 14100 13195
rect 13200 13150 14100 13155
rect -10550 13095 -9650 13100
rect -10550 13055 -10545 13095
rect -10505 13055 -10345 13095
rect -10305 13055 -10145 13095
rect -10105 13055 -9945 13095
rect -9905 13055 -9745 13095
rect -9705 13055 -9650 13095
rect -10550 13050 -9650 13055
rect 13200 13095 14100 13100
rect 13200 13055 13255 13095
rect 13295 13055 13655 13095
rect 13695 13055 14100 13095
rect 13200 13050 14100 13055
rect -10550 12995 -9650 13000
rect -10550 12955 -10545 12995
rect -10505 12955 -10345 12995
rect -10305 12955 -10145 12995
rect -10105 12955 -9945 12995
rect -9905 12955 -9745 12995
rect -9705 12955 -9650 12995
rect -10550 12950 -9650 12955
rect 13200 12995 14100 13000
rect 13200 12955 13255 12995
rect 13295 12955 13655 12995
rect 13695 12955 14100 12995
rect 13200 12950 14100 12955
rect 12600 12895 14000 12900
rect 12600 12855 13755 12895
rect 13795 12855 13955 12895
rect 13995 12855 14000 12895
rect 12600 12850 14000 12855
rect 12600 12795 13900 12800
rect 12600 12755 13855 12795
rect 13895 12755 13900 12795
rect 12600 12750 13900 12755
rect 12600 12695 14000 12700
rect 12600 12655 13755 12695
rect 13795 12655 13955 12695
rect 13995 12655 14000 12695
rect 12600 12650 14000 12655
rect -10550 12595 -9650 12600
rect -10550 12555 -10545 12595
rect -10505 12555 -10345 12595
rect -10305 12555 -10145 12595
rect -10105 12555 -9945 12595
rect -9905 12555 -9745 12595
rect -9705 12555 -9650 12595
rect -10550 12550 -9650 12555
rect 13200 12595 14100 12600
rect 13200 12555 13255 12595
rect 13295 12555 13655 12595
rect 13695 12555 14100 12595
rect 13200 12550 14100 12555
rect -10850 12295 -9650 12300
rect -10850 12255 -10845 12295
rect -10805 12255 -10795 12295
rect -10755 12255 -10745 12295
rect -10705 12255 -10695 12295
rect -10655 12255 -10645 12295
rect -10605 12255 -9650 12295
rect -10850 12250 -9650 12255
rect -10850 12195 -9650 12200
rect -10850 12155 -10845 12195
rect -10805 12155 -10795 12195
rect -10755 12155 -10745 12195
rect -10705 12155 -10695 12195
rect -10655 12155 -10645 12195
rect -10605 12155 -9650 12195
rect -10850 12150 -9650 12155
rect -10850 12095 -9650 12100
rect -10850 12055 -10845 12095
rect -10805 12055 -10795 12095
rect -10755 12055 -10745 12095
rect -10705 12055 -10695 12095
rect -10655 12055 -10645 12095
rect -10605 12055 -9650 12095
rect -10850 12050 -9650 12055
rect -10850 11995 -9650 12000
rect -10850 11955 -10845 11995
rect -10805 11955 -10795 11995
rect -10755 11955 -10745 11995
rect -10705 11955 -10695 11995
rect -10655 11955 -10645 11995
rect -10605 11955 -9650 11995
rect -10850 11950 -9650 11955
rect -10850 11895 -9650 11900
rect -10850 11855 -10845 11895
rect -10805 11855 -10795 11895
rect -10755 11855 -10745 11895
rect -10705 11855 -10695 11895
rect -10655 11855 -10645 11895
rect -10605 11855 -9650 11895
rect -10850 11850 -9650 11855
rect 13450 11895 14100 11900
rect 13450 11855 13455 11895
rect 13495 11855 14055 11895
rect 14095 11855 14100 11895
rect 13450 11850 14100 11855
rect -10850 11795 -9650 11800
rect -10850 11755 -10845 11795
rect -10805 11755 -10795 11795
rect -10755 11755 -10745 11795
rect -10705 11755 -10695 11795
rect -10655 11755 -10645 11795
rect -10605 11755 -9650 11795
rect -10850 11750 -9650 11755
rect 14150 11795 21850 15300
rect 14150 11755 14155 11795
rect 14195 11755 14205 11795
rect 14245 11755 14255 11795
rect 14295 11755 14305 11795
rect 14345 11755 14355 11795
rect 14395 11755 14405 11795
rect 14445 11755 14455 11795
rect 14495 11755 14505 11795
rect 14545 11755 14555 11795
rect 14595 11755 14605 11795
rect 14645 11755 14655 11795
rect 14695 11755 14705 11795
rect 14745 11755 14755 11795
rect 14795 11755 14805 11795
rect 14845 11755 14855 11795
rect 14895 11755 14905 11795
rect 14945 11755 14955 11795
rect 14995 11755 15005 11795
rect 15045 11755 15055 11795
rect 15095 11755 15105 11795
rect 15145 11755 15155 11795
rect 15195 11755 15205 11795
rect 15245 11755 15255 11795
rect 15295 11755 15305 11795
rect 15345 11755 15355 11795
rect 15395 11755 15405 11795
rect 15445 11755 15455 11795
rect 15495 11755 15505 11795
rect 15545 11755 15555 11795
rect 15595 11755 15605 11795
rect 15645 11755 15655 11795
rect 15695 11755 15705 11795
rect 15745 11755 15755 11795
rect 15795 11755 15805 11795
rect 15845 11755 15855 11795
rect 15895 11755 15905 11795
rect 15945 11755 15955 11795
rect 15995 11755 16005 11795
rect 16045 11755 16055 11795
rect 16095 11755 16105 11795
rect 16145 11755 16155 11795
rect 16195 11755 16205 11795
rect 16245 11755 16255 11795
rect 16295 11755 16305 11795
rect 16345 11755 16355 11795
rect 16395 11755 16405 11795
rect 16445 11755 16455 11795
rect 16495 11755 16505 11795
rect 16545 11755 16555 11795
rect 16595 11755 16605 11795
rect 16645 11755 16655 11795
rect 16695 11755 21705 11795
rect 21745 11755 21755 11795
rect 21795 11755 21805 11795
rect 21845 11755 21850 11795
rect 14150 11750 21850 11755
rect -10850 11695 -9650 11700
rect -10850 11655 -10845 11695
rect -10805 11655 -10795 11695
rect -10755 11655 -10745 11695
rect -10705 11655 -10695 11695
rect -10655 11655 -10645 11695
rect -10605 11655 -9650 11695
rect -10850 11650 -9650 11655
rect 13350 11695 21850 11700
rect 13350 11655 13355 11695
rect 13395 11655 13555 11695
rect 13595 11655 14155 11695
rect 14195 11655 14205 11695
rect 14245 11655 14255 11695
rect 14295 11655 14305 11695
rect 14345 11655 14355 11695
rect 14395 11655 14405 11695
rect 14445 11655 14455 11695
rect 14495 11655 14505 11695
rect 14545 11655 14555 11695
rect 14595 11655 14605 11695
rect 14645 11655 14655 11695
rect 14695 11655 14705 11695
rect 14745 11655 14755 11695
rect 14795 11655 14805 11695
rect 14845 11655 14855 11695
rect 14895 11655 14905 11695
rect 14945 11655 14955 11695
rect 14995 11655 15005 11695
rect 15045 11655 15055 11695
rect 15095 11655 15105 11695
rect 15145 11655 15155 11695
rect 15195 11655 15205 11695
rect 15245 11655 15255 11695
rect 15295 11655 15305 11695
rect 15345 11655 15355 11695
rect 15395 11655 15405 11695
rect 15445 11655 15455 11695
rect 15495 11655 15505 11695
rect 15545 11655 15555 11695
rect 15595 11655 15605 11695
rect 15645 11655 15655 11695
rect 15695 11655 15705 11695
rect 15745 11655 15755 11695
rect 15795 11655 15805 11695
rect 15845 11655 15855 11695
rect 15895 11655 15905 11695
rect 15945 11655 15955 11695
rect 15995 11655 16005 11695
rect 16045 11655 16055 11695
rect 16095 11655 16105 11695
rect 16145 11655 16155 11695
rect 16195 11655 16205 11695
rect 16245 11655 16255 11695
rect 16295 11655 16305 11695
rect 16345 11655 16355 11695
rect 16395 11655 16405 11695
rect 16445 11655 16455 11695
rect 16495 11655 16505 11695
rect 16545 11655 16555 11695
rect 16595 11655 16605 11695
rect 16645 11655 16655 11695
rect 16695 11655 21705 11695
rect 21745 11655 21755 11695
rect 21795 11655 21805 11695
rect 21845 11655 21850 11695
rect 13350 11650 21850 11655
rect -10950 11595 13200 11600
rect -10950 11555 -10945 11595
rect -10905 11590 13200 11595
rect -10905 11560 -9640 11590
rect -9610 11560 13200 11590
rect -10905 11555 13200 11560
rect -10950 11545 13200 11555
rect -10950 11505 -10945 11545
rect -10905 11540 13200 11545
rect -10905 11510 -9640 11540
rect -9610 11510 13200 11540
rect -10905 11505 13200 11510
rect -10950 11500 13200 11505
rect 13250 11595 13300 11600
rect 13250 11555 13255 11595
rect 13295 11555 13300 11595
rect 13250 11545 13300 11555
rect 13250 11505 13255 11545
rect 13295 11505 13300 11545
rect 13250 11500 13300 11505
rect 13650 11595 13700 11600
rect 13650 11555 13655 11595
rect 13695 11555 13700 11595
rect 13650 11545 13700 11555
rect 13650 11505 13655 11545
rect 13695 11505 13700 11545
rect 13650 11500 13700 11505
rect 14050 11595 21950 11600
rect 14050 11555 14055 11595
rect 14095 11555 21905 11595
rect 21945 11555 21950 11595
rect 14050 11545 21950 11555
rect 14050 11505 14055 11545
rect 14095 11505 21905 11545
rect 21945 11505 21950 11545
rect 14050 11500 21950 11505
rect -10850 11445 -9650 11450
rect -10850 11405 -10845 11445
rect -10805 11405 -10795 11445
rect -10755 11405 -10745 11445
rect -10705 11405 -10695 11445
rect -10655 11405 -10645 11445
rect -10605 11405 -9650 11445
rect -10850 11400 -9650 11405
rect 13750 11445 21850 11450
rect 13750 11405 13755 11445
rect 13795 11405 13955 11445
rect 13995 11405 14155 11445
rect 14195 11405 14205 11445
rect 14245 11405 14255 11445
rect 14295 11405 14305 11445
rect 14345 11405 14355 11445
rect 14395 11405 14405 11445
rect 14445 11405 14455 11445
rect 14495 11405 14505 11445
rect 14545 11405 14555 11445
rect 14595 11405 14605 11445
rect 14645 11405 14655 11445
rect 14695 11405 14705 11445
rect 14745 11405 14755 11445
rect 14795 11405 14805 11445
rect 14845 11405 14855 11445
rect 14895 11405 14905 11445
rect 14945 11405 14955 11445
rect 14995 11405 15005 11445
rect 15045 11405 15055 11445
rect 15095 11405 15105 11445
rect 15145 11405 15155 11445
rect 15195 11405 15205 11445
rect 15245 11405 15255 11445
rect 15295 11405 15305 11445
rect 15345 11405 15355 11445
rect 15395 11405 15405 11445
rect 15445 11405 15455 11445
rect 15495 11405 15505 11445
rect 15545 11405 15555 11445
rect 15595 11405 15605 11445
rect 15645 11405 15655 11445
rect 15695 11405 15705 11445
rect 15745 11405 15755 11445
rect 15795 11405 15805 11445
rect 15845 11405 15855 11445
rect 15895 11405 15905 11445
rect 15945 11405 15955 11445
rect 15995 11405 16005 11445
rect 16045 11405 16055 11445
rect 16095 11405 16105 11445
rect 16145 11405 16155 11445
rect 16195 11405 16205 11445
rect 16245 11405 16255 11445
rect 16295 11405 16305 11445
rect 16345 11405 16355 11445
rect 16395 11405 16405 11445
rect 16445 11405 16455 11445
rect 16495 11405 16505 11445
rect 16545 11405 16555 11445
rect 16595 11405 16605 11445
rect 16645 11405 16655 11445
rect 16695 11405 21705 11445
rect 21745 11405 21755 11445
rect 21795 11405 21805 11445
rect 21845 11405 21850 11445
rect 13750 11400 21850 11405
rect -10850 11345 -9650 11350
rect -10850 11305 -10845 11345
rect -10805 11305 -10795 11345
rect -10755 11305 -10745 11345
rect -10705 11305 -10695 11345
rect -10655 11305 -10645 11345
rect -10605 11305 -9650 11345
rect -10850 11300 -9650 11305
rect 14150 11345 21850 11350
rect 14150 11305 14155 11345
rect 14195 11305 14205 11345
rect 14245 11305 14255 11345
rect 14295 11305 14305 11345
rect 14345 11305 14355 11345
rect 14395 11305 14405 11345
rect 14445 11305 14455 11345
rect 14495 11305 14505 11345
rect 14545 11305 14555 11345
rect 14595 11305 14605 11345
rect 14645 11305 14655 11345
rect 14695 11305 14705 11345
rect 14745 11305 14755 11345
rect 14795 11305 14805 11345
rect 14845 11305 14855 11345
rect 14895 11305 14905 11345
rect 14945 11305 14955 11345
rect 14995 11305 15005 11345
rect 15045 11305 15055 11345
rect 15095 11305 15105 11345
rect 15145 11305 15155 11345
rect 15195 11305 15205 11345
rect 15245 11305 15255 11345
rect 15295 11305 15305 11345
rect 15345 11305 15355 11345
rect 15395 11305 15405 11345
rect 15445 11305 15455 11345
rect 15495 11305 15505 11345
rect 15545 11305 15555 11345
rect 15595 11305 15605 11345
rect 15645 11305 15655 11345
rect 15695 11305 15705 11345
rect 15745 11305 15755 11345
rect 15795 11305 15805 11345
rect 15845 11305 15855 11345
rect 15895 11305 15905 11345
rect 15945 11305 15955 11345
rect 15995 11305 16005 11345
rect 16045 11305 16055 11345
rect 16095 11305 16105 11345
rect 16145 11305 16155 11345
rect 16195 11305 16205 11345
rect 16245 11305 16255 11345
rect 16295 11305 16305 11345
rect 16345 11305 16355 11345
rect 16395 11305 16405 11345
rect 16445 11305 16455 11345
rect 16495 11305 16505 11345
rect 16545 11305 16555 11345
rect 16595 11305 16605 11345
rect 16645 11305 16655 11345
rect 16695 11305 21705 11345
rect 21745 11305 21755 11345
rect 21795 11305 21805 11345
rect 21845 11305 21850 11345
rect -10850 11245 -9650 11250
rect -10850 11205 -10845 11245
rect -10805 11205 -10795 11245
rect -10755 11205 -10745 11245
rect -10705 11205 -10695 11245
rect -10655 11205 -10645 11245
rect -10605 11205 -9650 11245
rect -10850 11200 -9650 11205
rect 13850 11245 14100 11250
rect 13850 11205 13855 11245
rect 13895 11205 14055 11245
rect 14095 11205 14100 11245
rect 13850 11200 14100 11205
rect -10850 11145 -9650 11150
rect -10850 11105 -10845 11145
rect -10805 11105 -10795 11145
rect -10755 11105 -10745 11145
rect -10705 11105 -10695 11145
rect -10655 11105 -10645 11145
rect -10605 11105 -9650 11145
rect -10850 11100 -9650 11105
rect -10850 11045 -9650 11050
rect -10850 11005 -10845 11045
rect -10805 11005 -10795 11045
rect -10755 11005 -10745 11045
rect -10705 11005 -10695 11045
rect -10655 11005 -10645 11045
rect -10605 11005 -9650 11045
rect -10850 11000 -9650 11005
rect -10850 10945 -9650 10950
rect -10850 10905 -10845 10945
rect -10805 10905 -10795 10945
rect -10755 10905 -10745 10945
rect -10705 10905 -10695 10945
rect -10655 10905 -10645 10945
rect -10605 10905 -9650 10945
rect -10850 10900 -9650 10905
rect -10850 10845 -9650 10850
rect -10850 10805 -10845 10845
rect -10805 10805 -10795 10845
rect -10755 10805 -10745 10845
rect -10705 10805 -10695 10845
rect -10655 10805 -10645 10845
rect -10605 10805 -9650 10845
rect -10850 10800 -9650 10805
rect -10550 10545 -9650 10550
rect -10550 10505 -10545 10545
rect -10505 10505 -10345 10545
rect -10305 10505 -10145 10545
rect -10105 10505 -9945 10545
rect -9905 10505 -9745 10545
rect -9705 10505 -9650 10545
rect -10550 10500 -9650 10505
rect 13200 10545 14100 10550
rect 13200 10505 13255 10545
rect 13295 10505 13655 10545
rect 13695 10505 14100 10545
rect 13200 10500 14100 10505
rect 12600 10445 14000 10450
rect 12600 10405 13755 10445
rect 13795 10405 13955 10445
rect 13995 10405 14000 10445
rect 12600 10400 14000 10405
rect 12600 10345 13900 10350
rect 12600 10305 13855 10345
rect 13895 10305 13900 10345
rect 12600 10300 13900 10305
rect 12600 10245 14000 10250
rect 12600 10205 13755 10245
rect 13795 10205 13955 10245
rect 13995 10205 14000 10245
rect 12600 10200 14000 10205
rect -10550 10145 -9650 10150
rect -10550 10105 -10545 10145
rect -10505 10105 -10345 10145
rect -10305 10105 -10145 10145
rect -10105 10105 -9945 10145
rect -9905 10105 -9745 10145
rect -9705 10105 -9650 10145
rect -10550 10100 -9650 10105
rect 13200 10145 14100 10150
rect 13200 10105 13255 10145
rect 13295 10105 13655 10145
rect 13695 10105 14100 10145
rect 13200 10100 14100 10105
rect -10550 10045 -9650 10050
rect -10550 10005 -10545 10045
rect -10505 10005 -10345 10045
rect -10305 10005 -10145 10045
rect -10105 10005 -9945 10045
rect -9905 10005 -9745 10045
rect -9705 10005 -9650 10045
rect -10550 10000 -9650 10005
rect 13200 10045 14100 10050
rect 13200 10005 13255 10045
rect 13295 10005 13655 10045
rect 13695 10005 14100 10045
rect 13200 10000 14100 10005
rect -10550 9945 -9650 9950
rect -10550 9905 -10545 9945
rect -10505 9905 -10345 9945
rect -10305 9905 -10145 9945
rect -10105 9905 -9945 9945
rect -9905 9905 -9745 9945
rect -9705 9905 -9650 9945
rect -10550 9900 -9650 9905
rect 13200 9945 14100 9950
rect 13200 9905 13255 9945
rect 13295 9905 13655 9945
rect 13695 9905 14100 9945
rect 13200 9900 14100 9905
rect -10050 9845 -9050 9850
rect -10050 9805 -10045 9845
rect -10005 9805 -9050 9845
rect -10050 9800 -9050 9805
rect 13200 9845 14100 9850
rect 13200 9805 13255 9845
rect 13295 9805 13655 9845
rect 13695 9805 14100 9845
rect 13200 9800 14100 9805
rect -10550 9745 -9650 9750
rect -10550 9705 -10545 9745
rect -10505 9705 -10345 9745
rect -10305 9705 -10145 9745
rect -10105 9705 -9945 9745
rect -9905 9705 -9745 9745
rect -9705 9705 -9650 9745
rect -10550 9700 -9650 9705
rect 13200 9745 14100 9750
rect 13200 9705 13255 9745
rect 13295 9705 13655 9745
rect 13695 9705 14100 9745
rect 13200 9700 14100 9705
rect -9500 9645 -9450 9650
rect -9500 9605 -9495 9645
rect -9455 9605 -9450 9645
rect -9500 9600 -9450 9605
rect -9350 9645 -9300 9650
rect -9350 9605 -9345 9645
rect -9305 9605 -9300 9645
rect -9350 9600 -9300 9605
rect -10550 9545 -9650 9550
rect -10550 9505 -10545 9545
rect -10505 9505 -10345 9545
rect -10305 9505 -10145 9545
rect -10105 9505 -9945 9545
rect -9905 9505 -9745 9545
rect -9705 9505 -9650 9545
rect -10550 9500 -9650 9505
rect 13200 9545 14100 9550
rect 13200 9505 13255 9545
rect 13295 9505 13655 9545
rect 13695 9505 14100 9545
rect 13200 9500 14100 9505
rect -9850 9445 -9050 9450
rect -9850 9405 -9845 9445
rect -9805 9405 -9050 9445
rect -9850 9400 -9050 9405
rect 13200 9445 14100 9450
rect 13200 9405 13255 9445
rect 13295 9405 13655 9445
rect 13695 9405 14100 9445
rect 13200 9400 14100 9405
rect -10550 9345 -9650 9350
rect -10550 9305 -10545 9345
rect -10505 9305 -10345 9345
rect -10305 9305 -10145 9345
rect -10105 9305 -9945 9345
rect -9905 9305 -9745 9345
rect -9705 9305 -9650 9345
rect -10550 9300 -9650 9305
rect 13200 9345 14100 9350
rect 13200 9305 13255 9345
rect 13295 9305 13655 9345
rect 13695 9305 14100 9345
rect 13200 9300 14100 9305
rect -10550 9245 -9650 9250
rect -10550 9205 -10545 9245
rect -10505 9205 -10345 9245
rect -10305 9205 -10145 9245
rect -10105 9205 -9945 9245
rect -9905 9205 -9745 9245
rect -9705 9205 -9650 9245
rect -10550 9200 -9650 9205
rect 13200 9245 14100 9250
rect 13200 9205 13255 9245
rect 13295 9205 13655 9245
rect 13695 9205 14100 9245
rect 13200 9200 14100 9205
rect -10550 9145 -9650 9150
rect -10550 9105 -10545 9145
rect -10505 9105 -10345 9145
rect -10305 9105 -10145 9145
rect -10105 9105 -9945 9145
rect -9905 9105 -9745 9145
rect -9705 9105 -9650 9145
rect -10550 9100 -9650 9105
rect 13200 9145 14100 9150
rect 13200 9105 13255 9145
rect 13295 9105 13655 9145
rect 13695 9105 14100 9145
rect 13200 9100 14100 9105
rect 12600 9045 13600 9050
rect 12600 9005 13355 9045
rect 13395 9005 13555 9045
rect 13595 9005 13600 9045
rect 12600 9000 13600 9005
rect 12600 8945 13500 8950
rect 12600 8905 13455 8945
rect 13495 8905 13500 8945
rect 12600 8900 13500 8905
rect 12600 8845 13600 8850
rect 12600 8805 13355 8845
rect 13395 8805 13555 8845
rect 13595 8805 13600 8845
rect 12600 8800 13600 8805
rect -10550 8745 -9650 8750
rect -10550 8705 -10545 8745
rect -10505 8705 -10345 8745
rect -10305 8705 -10145 8745
rect -10105 8705 -9945 8745
rect -9905 8705 -9745 8745
rect -9705 8705 -9650 8745
rect -10550 8700 -9650 8705
rect 13200 8745 14100 8750
rect 13200 8705 13255 8745
rect 13295 8705 13655 8745
rect 13695 8705 14055 8745
rect 14095 8705 14100 8745
rect 13200 8700 14100 8705
rect -10850 8445 -9650 8450
rect -10850 8405 -10845 8445
rect -10805 8405 -10795 8445
rect -10755 8405 -10745 8445
rect -10705 8405 -10695 8445
rect -10655 8405 -10645 8445
rect -10605 8405 -9650 8445
rect -10850 8400 -9650 8405
rect -10850 8345 -9650 8350
rect -10850 8305 -10845 8345
rect -10805 8305 -10795 8345
rect -10755 8305 -10745 8345
rect -10705 8305 -10695 8345
rect -10655 8305 -10645 8345
rect -10605 8305 -9650 8345
rect -10850 8300 -9650 8305
rect -10850 8245 -9650 8250
rect -10850 8205 -10845 8245
rect -10805 8205 -10795 8245
rect -10755 8205 -10745 8245
rect -10705 8205 -10695 8245
rect -10655 8205 -10645 8245
rect -10605 8205 -9650 8245
rect -10850 8200 -9650 8205
rect -10850 8145 -9650 8150
rect -10850 8105 -10845 8145
rect -10805 8105 -10795 8145
rect -10755 8105 -10745 8145
rect -10705 8105 -10695 8145
rect -10655 8105 -10645 8145
rect -10605 8105 -9650 8145
rect -10850 8100 -9650 8105
rect -10850 8045 -9650 8050
rect -10850 8005 -10845 8045
rect -10805 8005 -10795 8045
rect -10755 8005 -10745 8045
rect -10705 8005 -10695 8045
rect -10655 8005 -10645 8045
rect -10605 8005 -9650 8045
rect -10850 8000 -9650 8005
rect -10850 7945 -9650 7950
rect -10850 7905 -10845 7945
rect -10805 7905 -10795 7945
rect -10755 7905 -10745 7945
rect -10705 7905 -10695 7945
rect -10655 7905 -10645 7945
rect -10605 7905 -9650 7945
rect -10850 7900 -9650 7905
rect -10850 7845 -9650 7850
rect -10850 7805 -10845 7845
rect -10805 7805 -10795 7845
rect -10755 7805 -10745 7845
rect -10705 7805 -10695 7845
rect -10655 7805 -10645 7845
rect -10605 7805 -9650 7845
rect -10850 7800 -9650 7805
rect 14150 7800 21850 11305
rect 13250 7745 21950 7750
rect 13250 7705 13255 7745
rect 13295 7705 13655 7745
rect 13695 7705 21905 7745
rect 21945 7705 21950 7745
rect 13250 7700 21950 7705
<< via3 >>
rect 14055 15355 14095 15395
rect 21905 15355 21945 15395
rect -10845 15255 -10805 15295
rect -10795 15255 -10755 15295
rect -10745 15255 -10705 15295
rect -10695 15255 -10655 15295
rect -10645 15255 -10605 15295
rect -10845 15155 -10805 15195
rect -10795 15155 -10755 15195
rect -10745 15155 -10705 15195
rect -10695 15155 -10655 15195
rect -10645 15155 -10605 15195
rect -10845 15055 -10805 15095
rect -10795 15055 -10755 15095
rect -10745 15055 -10705 15095
rect -10695 15055 -10655 15095
rect -10645 15055 -10605 15095
rect -10845 14955 -10805 14995
rect -10795 14955 -10755 14995
rect -10745 14955 -10705 14995
rect -10695 14955 -10655 14995
rect -10645 14955 -10605 14995
rect -10845 14855 -10805 14895
rect -10795 14855 -10755 14895
rect -10745 14855 -10705 14895
rect -10695 14855 -10655 14895
rect -10645 14855 -10605 14895
rect -10845 14755 -10805 14795
rect -10795 14755 -10755 14795
rect -10745 14755 -10705 14795
rect -10695 14755 -10655 14795
rect -10645 14755 -10605 14795
rect -10845 14655 -10805 14695
rect -10795 14655 -10755 14695
rect -10745 14655 -10705 14695
rect -10695 14655 -10655 14695
rect -10645 14655 -10605 14695
rect -10545 14355 -10505 14395
rect -10345 14355 -10305 14395
rect -10145 14355 -10105 14395
rect -9945 14355 -9905 14395
rect -9745 14355 -9705 14395
rect 13255 14355 13295 14395
rect 13655 14355 13695 14395
rect 13355 14255 13395 14295
rect 13555 14255 13595 14295
rect 13455 14155 13495 14195
rect 13355 14055 13395 14095
rect 13555 14055 13595 14095
rect -10545 13955 -10505 13995
rect -10345 13955 -10305 13995
rect -10145 13955 -10105 13995
rect -9945 13955 -9905 13995
rect -9745 13955 -9705 13995
rect 13255 13955 13295 13995
rect 13655 13955 13695 13995
rect -10545 13855 -10505 13895
rect -10345 13855 -10305 13895
rect -10145 13855 -10105 13895
rect -9945 13855 -9905 13895
rect -9745 13855 -9705 13895
rect 13255 13855 13295 13895
rect 13655 13855 13695 13895
rect -10545 13755 -10505 13795
rect -10345 13755 -10305 13795
rect -10145 13755 -10105 13795
rect -9945 13755 -9905 13795
rect -9745 13755 -9705 13795
rect 13255 13755 13295 13795
rect 13655 13755 13695 13795
rect -10245 13655 -10205 13695
rect 13255 13655 13295 13695
rect 13655 13655 13695 13695
rect -10545 13555 -10505 13595
rect -10345 13555 -10305 13595
rect -10145 13555 -10105 13595
rect -9945 13555 -9905 13595
rect -9745 13555 -9705 13595
rect 13255 13555 13295 13595
rect 13655 13555 13695 13595
rect -9495 13490 -9455 13495
rect -9495 13460 -9490 13490
rect -9490 13460 -9460 13490
rect -9460 13460 -9455 13490
rect -9495 13455 -9455 13460
rect -9345 13490 -9305 13495
rect -9345 13460 -9340 13490
rect -9340 13460 -9310 13490
rect -9310 13460 -9305 13490
rect -9345 13455 -9305 13460
rect -10545 13355 -10505 13395
rect -10345 13355 -10305 13395
rect -10145 13355 -10105 13395
rect -9945 13355 -9905 13395
rect -9745 13355 -9705 13395
rect 13255 13355 13295 13395
rect 13655 13355 13695 13395
rect -10445 13255 -10405 13295
rect 13255 13255 13295 13295
rect 13655 13255 13695 13295
rect -10545 13155 -10505 13195
rect -10345 13155 -10305 13195
rect -10145 13155 -10105 13195
rect -9945 13155 -9905 13195
rect -9745 13155 -9705 13195
rect 13255 13155 13295 13195
rect 13655 13155 13695 13195
rect -10545 13055 -10505 13095
rect -10345 13055 -10305 13095
rect -10145 13055 -10105 13095
rect -9945 13055 -9905 13095
rect -9745 13055 -9705 13095
rect 13255 13055 13295 13095
rect 13655 13055 13695 13095
rect -10545 12955 -10505 12995
rect -10345 12955 -10305 12995
rect -10145 12955 -10105 12995
rect -9945 12955 -9905 12995
rect -9745 12955 -9705 12995
rect 13255 12955 13295 12995
rect 13655 12955 13695 12995
rect 13755 12855 13795 12895
rect 13955 12855 13995 12895
rect 13855 12755 13895 12795
rect 13755 12655 13795 12695
rect 13955 12655 13995 12695
rect -10545 12555 -10505 12595
rect -10345 12555 -10305 12595
rect -10145 12555 -10105 12595
rect -9945 12555 -9905 12595
rect -9745 12555 -9705 12595
rect 13255 12555 13295 12595
rect 13655 12555 13695 12595
rect -10845 12255 -10805 12295
rect -10795 12255 -10755 12295
rect -10745 12255 -10705 12295
rect -10695 12255 -10655 12295
rect -10645 12255 -10605 12295
rect -10845 12155 -10805 12195
rect -10795 12155 -10755 12195
rect -10745 12155 -10705 12195
rect -10695 12155 -10655 12195
rect -10645 12155 -10605 12195
rect -10845 12055 -10805 12095
rect -10795 12055 -10755 12095
rect -10745 12055 -10705 12095
rect -10695 12055 -10655 12095
rect -10645 12055 -10605 12095
rect -10845 11955 -10805 11995
rect -10795 11955 -10755 11995
rect -10745 11955 -10705 11995
rect -10695 11955 -10655 11995
rect -10645 11955 -10605 11995
rect -10845 11855 -10805 11895
rect -10795 11855 -10755 11895
rect -10745 11855 -10705 11895
rect -10695 11855 -10655 11895
rect -10645 11855 -10605 11895
rect 13455 11855 13495 11895
rect 14055 11855 14095 11895
rect -10845 11755 -10805 11795
rect -10795 11755 -10755 11795
rect -10745 11755 -10705 11795
rect -10695 11755 -10655 11795
rect -10645 11755 -10605 11795
rect 14155 11755 14195 11795
rect 14205 11755 14245 11795
rect 14255 11755 14295 11795
rect 14305 11755 14345 11795
rect 14355 11755 14395 11795
rect 14405 11755 14445 11795
rect 14455 11755 14495 11795
rect 14505 11755 14545 11795
rect 14555 11755 14595 11795
rect 14605 11755 14645 11795
rect 14655 11755 14695 11795
rect 14705 11755 14745 11795
rect 14755 11755 14795 11795
rect 14805 11755 14845 11795
rect 14855 11755 14895 11795
rect 14905 11755 14945 11795
rect 14955 11755 14995 11795
rect 15005 11755 15045 11795
rect 15055 11755 15095 11795
rect 15105 11755 15145 11795
rect 15155 11755 15195 11795
rect 15205 11755 15245 11795
rect 15255 11755 15295 11795
rect 15305 11755 15345 11795
rect 15355 11755 15395 11795
rect 15405 11755 15445 11795
rect 15455 11755 15495 11795
rect 15505 11755 15545 11795
rect 15555 11755 15595 11795
rect 15605 11755 15645 11795
rect 15655 11755 15695 11795
rect 15705 11755 15745 11795
rect 15755 11755 15795 11795
rect 15805 11755 15845 11795
rect 15855 11755 15895 11795
rect 15905 11755 15945 11795
rect 15955 11755 15995 11795
rect 16005 11755 16045 11795
rect 16055 11755 16095 11795
rect 16105 11755 16145 11795
rect 16155 11755 16195 11795
rect 16205 11755 16245 11795
rect 16255 11755 16295 11795
rect 16305 11755 16345 11795
rect 16355 11755 16395 11795
rect 16405 11755 16445 11795
rect 16455 11755 16495 11795
rect 16505 11755 16545 11795
rect 16555 11755 16595 11795
rect 16605 11755 16645 11795
rect 16655 11755 16695 11795
rect 21705 11755 21745 11795
rect 21755 11755 21795 11795
rect 21805 11755 21845 11795
rect -10845 11655 -10805 11695
rect -10795 11655 -10755 11695
rect -10745 11655 -10705 11695
rect -10695 11655 -10655 11695
rect -10645 11655 -10605 11695
rect 13355 11655 13395 11695
rect 13555 11655 13595 11695
rect 14155 11655 14195 11695
rect 14205 11655 14245 11695
rect 14255 11655 14295 11695
rect 14305 11655 14345 11695
rect 14355 11655 14395 11695
rect 14405 11655 14445 11695
rect 14455 11655 14495 11695
rect 14505 11655 14545 11695
rect 14555 11655 14595 11695
rect 14605 11655 14645 11695
rect 14655 11655 14695 11695
rect 14705 11655 14745 11695
rect 14755 11655 14795 11695
rect 14805 11655 14845 11695
rect 14855 11655 14895 11695
rect 14905 11655 14945 11695
rect 14955 11655 14995 11695
rect 15005 11655 15045 11695
rect 15055 11655 15095 11695
rect 15105 11655 15145 11695
rect 15155 11655 15195 11695
rect 15205 11655 15245 11695
rect 15255 11655 15295 11695
rect 15305 11655 15345 11695
rect 15355 11655 15395 11695
rect 15405 11655 15445 11695
rect 15455 11655 15495 11695
rect 15505 11655 15545 11695
rect 15555 11655 15595 11695
rect 15605 11655 15645 11695
rect 15655 11655 15695 11695
rect 15705 11655 15745 11695
rect 15755 11655 15795 11695
rect 15805 11655 15845 11695
rect 15855 11655 15895 11695
rect 15905 11655 15945 11695
rect 15955 11655 15995 11695
rect 16005 11655 16045 11695
rect 16055 11655 16095 11695
rect 16105 11655 16145 11695
rect 16155 11655 16195 11695
rect 16205 11655 16245 11695
rect 16255 11655 16295 11695
rect 16305 11655 16345 11695
rect 16355 11655 16395 11695
rect 16405 11655 16445 11695
rect 16455 11655 16495 11695
rect 16505 11655 16545 11695
rect 16555 11655 16595 11695
rect 16605 11655 16645 11695
rect 16655 11655 16695 11695
rect 21705 11655 21745 11695
rect 21755 11655 21795 11695
rect 21805 11655 21845 11695
rect -10945 11590 -10905 11595
rect -10945 11560 -10940 11590
rect -10940 11560 -10910 11590
rect -10910 11560 -10905 11590
rect -10945 11555 -10905 11560
rect -10945 11540 -10905 11545
rect -10945 11510 -10940 11540
rect -10940 11510 -10910 11540
rect -10910 11510 -10905 11540
rect -10945 11505 -10905 11510
rect 13255 11555 13295 11595
rect 13255 11505 13295 11545
rect 13655 11555 13695 11595
rect 13655 11505 13695 11545
rect 14055 11555 14095 11595
rect 21905 11555 21945 11595
rect 14055 11505 14095 11545
rect 21905 11505 21945 11545
rect -10845 11405 -10805 11445
rect -10795 11405 -10755 11445
rect -10745 11405 -10705 11445
rect -10695 11405 -10655 11445
rect -10645 11405 -10605 11445
rect 13755 11405 13795 11445
rect 13955 11405 13995 11445
rect 14155 11405 14195 11445
rect 14205 11405 14245 11445
rect 14255 11405 14295 11445
rect 14305 11405 14345 11445
rect 14355 11405 14395 11445
rect 14405 11405 14445 11445
rect 14455 11405 14495 11445
rect 14505 11405 14545 11445
rect 14555 11405 14595 11445
rect 14605 11405 14645 11445
rect 14655 11405 14695 11445
rect 14705 11405 14745 11445
rect 14755 11405 14795 11445
rect 14805 11405 14845 11445
rect 14855 11405 14895 11445
rect 14905 11405 14945 11445
rect 14955 11405 14995 11445
rect 15005 11405 15045 11445
rect 15055 11405 15095 11445
rect 15105 11405 15145 11445
rect 15155 11405 15195 11445
rect 15205 11405 15245 11445
rect 15255 11405 15295 11445
rect 15305 11405 15345 11445
rect 15355 11405 15395 11445
rect 15405 11405 15445 11445
rect 15455 11405 15495 11445
rect 15505 11405 15545 11445
rect 15555 11405 15595 11445
rect 15605 11405 15645 11445
rect 15655 11405 15695 11445
rect 15705 11405 15745 11445
rect 15755 11405 15795 11445
rect 15805 11405 15845 11445
rect 15855 11405 15895 11445
rect 15905 11405 15945 11445
rect 15955 11405 15995 11445
rect 16005 11405 16045 11445
rect 16055 11405 16095 11445
rect 16105 11405 16145 11445
rect 16155 11405 16195 11445
rect 16205 11405 16245 11445
rect 16255 11405 16295 11445
rect 16305 11405 16345 11445
rect 16355 11405 16395 11445
rect 16405 11405 16445 11445
rect 16455 11405 16495 11445
rect 16505 11405 16545 11445
rect 16555 11405 16595 11445
rect 16605 11405 16645 11445
rect 16655 11405 16695 11445
rect 21705 11405 21745 11445
rect 21755 11405 21795 11445
rect 21805 11405 21845 11445
rect -10845 11305 -10805 11345
rect -10795 11305 -10755 11345
rect -10745 11305 -10705 11345
rect -10695 11305 -10655 11345
rect -10645 11305 -10605 11345
rect 14155 11305 14195 11345
rect 14205 11305 14245 11345
rect 14255 11305 14295 11345
rect 14305 11305 14345 11345
rect 14355 11305 14395 11345
rect 14405 11305 14445 11345
rect 14455 11305 14495 11345
rect 14505 11305 14545 11345
rect 14555 11305 14595 11345
rect 14605 11305 14645 11345
rect 14655 11305 14695 11345
rect 14705 11305 14745 11345
rect 14755 11305 14795 11345
rect 14805 11305 14845 11345
rect 14855 11305 14895 11345
rect 14905 11305 14945 11345
rect 14955 11305 14995 11345
rect 15005 11305 15045 11345
rect 15055 11305 15095 11345
rect 15105 11305 15145 11345
rect 15155 11305 15195 11345
rect 15205 11305 15245 11345
rect 15255 11305 15295 11345
rect 15305 11305 15345 11345
rect 15355 11305 15395 11345
rect 15405 11305 15445 11345
rect 15455 11305 15495 11345
rect 15505 11305 15545 11345
rect 15555 11305 15595 11345
rect 15605 11305 15645 11345
rect 15655 11305 15695 11345
rect 15705 11305 15745 11345
rect 15755 11305 15795 11345
rect 15805 11305 15845 11345
rect 15855 11305 15895 11345
rect 15905 11305 15945 11345
rect 15955 11305 15995 11345
rect 16005 11305 16045 11345
rect 16055 11305 16095 11345
rect 16105 11305 16145 11345
rect 16155 11305 16195 11345
rect 16205 11305 16245 11345
rect 16255 11305 16295 11345
rect 16305 11305 16345 11345
rect 16355 11305 16395 11345
rect 16405 11305 16445 11345
rect 16455 11305 16495 11345
rect 16505 11305 16545 11345
rect 16555 11305 16595 11345
rect 16605 11305 16645 11345
rect 16655 11305 16695 11345
rect 21705 11305 21745 11345
rect 21755 11305 21795 11345
rect 21805 11305 21845 11345
rect -10845 11205 -10805 11245
rect -10795 11205 -10755 11245
rect -10745 11205 -10705 11245
rect -10695 11205 -10655 11245
rect -10645 11205 -10605 11245
rect 13855 11205 13895 11245
rect 14055 11205 14095 11245
rect -10845 11105 -10805 11145
rect -10795 11105 -10755 11145
rect -10745 11105 -10705 11145
rect -10695 11105 -10655 11145
rect -10645 11105 -10605 11145
rect -10845 11005 -10805 11045
rect -10795 11005 -10755 11045
rect -10745 11005 -10705 11045
rect -10695 11005 -10655 11045
rect -10645 11005 -10605 11045
rect -10845 10905 -10805 10945
rect -10795 10905 -10755 10945
rect -10745 10905 -10705 10945
rect -10695 10905 -10655 10945
rect -10645 10905 -10605 10945
rect -10845 10805 -10805 10845
rect -10795 10805 -10755 10845
rect -10745 10805 -10705 10845
rect -10695 10805 -10655 10845
rect -10645 10805 -10605 10845
rect -10545 10505 -10505 10545
rect -10345 10505 -10305 10545
rect -10145 10505 -10105 10545
rect -9945 10505 -9905 10545
rect -9745 10505 -9705 10545
rect 13255 10505 13295 10545
rect 13655 10505 13695 10545
rect 13755 10405 13795 10445
rect 13955 10405 13995 10445
rect 13855 10305 13895 10345
rect 13755 10205 13795 10245
rect 13955 10205 13995 10245
rect -10545 10105 -10505 10145
rect -10345 10105 -10305 10145
rect -10145 10105 -10105 10145
rect -9945 10105 -9905 10145
rect -9745 10105 -9705 10145
rect 13255 10105 13295 10145
rect 13655 10105 13695 10145
rect -10545 10005 -10505 10045
rect -10345 10005 -10305 10045
rect -10145 10005 -10105 10045
rect -9945 10005 -9905 10045
rect -9745 10005 -9705 10045
rect 13255 10005 13295 10045
rect 13655 10005 13695 10045
rect -10545 9905 -10505 9945
rect -10345 9905 -10305 9945
rect -10145 9905 -10105 9945
rect -9945 9905 -9905 9945
rect -9745 9905 -9705 9945
rect 13255 9905 13295 9945
rect 13655 9905 13695 9945
rect -10045 9805 -10005 9845
rect 13255 9805 13295 9845
rect 13655 9805 13695 9845
rect -10545 9705 -10505 9745
rect -10345 9705 -10305 9745
rect -10145 9705 -10105 9745
rect -9945 9705 -9905 9745
rect -9745 9705 -9705 9745
rect 13255 9705 13295 9745
rect 13655 9705 13695 9745
rect -9495 9640 -9455 9645
rect -9495 9610 -9490 9640
rect -9490 9610 -9460 9640
rect -9460 9610 -9455 9640
rect -9495 9605 -9455 9610
rect -9345 9640 -9305 9645
rect -9345 9610 -9340 9640
rect -9340 9610 -9310 9640
rect -9310 9610 -9305 9640
rect -9345 9605 -9305 9610
rect -10545 9505 -10505 9545
rect -10345 9505 -10305 9545
rect -10145 9505 -10105 9545
rect -9945 9505 -9905 9545
rect -9745 9505 -9705 9545
rect 13255 9505 13295 9545
rect 13655 9505 13695 9545
rect -9845 9405 -9805 9445
rect 13255 9405 13295 9445
rect 13655 9405 13695 9445
rect -10545 9305 -10505 9345
rect -10345 9305 -10305 9345
rect -10145 9305 -10105 9345
rect -9945 9305 -9905 9345
rect -9745 9305 -9705 9345
rect 13255 9305 13295 9345
rect 13655 9305 13695 9345
rect -10545 9205 -10505 9245
rect -10345 9205 -10305 9245
rect -10145 9205 -10105 9245
rect -9945 9205 -9905 9245
rect -9745 9205 -9705 9245
rect 13255 9205 13295 9245
rect 13655 9205 13695 9245
rect -10545 9105 -10505 9145
rect -10345 9105 -10305 9145
rect -10145 9105 -10105 9145
rect -9945 9105 -9905 9145
rect -9745 9105 -9705 9145
rect 13255 9105 13295 9145
rect 13655 9105 13695 9145
rect 13355 9005 13395 9045
rect 13555 9005 13595 9045
rect 13455 8905 13495 8945
rect 13355 8805 13395 8845
rect 13555 8805 13595 8845
rect -10545 8705 -10505 8745
rect -10345 8705 -10305 8745
rect -10145 8705 -10105 8745
rect -9945 8705 -9905 8745
rect -9745 8705 -9705 8745
rect 13255 8705 13295 8745
rect 13655 8705 13695 8745
rect 14055 8705 14095 8745
rect -10845 8405 -10805 8445
rect -10795 8405 -10755 8445
rect -10745 8405 -10705 8445
rect -10695 8405 -10655 8445
rect -10645 8405 -10605 8445
rect -10845 8305 -10805 8345
rect -10795 8305 -10755 8345
rect -10745 8305 -10705 8345
rect -10695 8305 -10655 8345
rect -10645 8305 -10605 8345
rect -10845 8205 -10805 8245
rect -10795 8205 -10755 8245
rect -10745 8205 -10705 8245
rect -10695 8205 -10655 8245
rect -10645 8205 -10605 8245
rect -10845 8105 -10805 8145
rect -10795 8105 -10755 8145
rect -10745 8105 -10705 8145
rect -10695 8105 -10655 8145
rect -10645 8105 -10605 8145
rect -10845 8005 -10805 8045
rect -10795 8005 -10755 8045
rect -10745 8005 -10705 8045
rect -10695 8005 -10655 8045
rect -10645 8005 -10605 8045
rect -10845 7905 -10805 7945
rect -10795 7905 -10755 7945
rect -10745 7905 -10705 7945
rect -10695 7905 -10655 7945
rect -10645 7905 -10605 7945
rect -10845 7805 -10805 7845
rect -10795 7805 -10755 7845
rect -10745 7805 -10705 7845
rect -10695 7805 -10655 7845
rect -10645 7805 -10605 7845
rect 13255 7705 13295 7745
rect 13655 7705 13695 7745
rect 21905 7705 21945 7745
<< mimcap >>
rect 14200 15200 21800 15250
rect 14200 11950 14250 15200
rect 21750 11950 21800 15200
rect 14200 11900 21800 11950
rect 14200 11150 21800 11200
rect 14200 7900 14250 11150
rect 21750 7900 21800 11150
rect 14200 7850 21800 7900
<< mimcapcontact >>
rect 14250 11950 21750 15200
rect 14250 7900 21750 11150
<< metal4 >>
rect -10950 11595 -10900 15400
rect -10950 11555 -10945 11595
rect -10905 11555 -10900 11595
rect -10950 11545 -10900 11555
rect -10950 11505 -10945 11545
rect -10905 11505 -10900 11545
rect -10950 7700 -10900 11505
rect -10850 15295 -10600 15400
rect -10850 15255 -10845 15295
rect -10805 15255 -10795 15295
rect -10755 15255 -10745 15295
rect -10705 15255 -10695 15295
rect -10655 15255 -10645 15295
rect -10605 15255 -10600 15295
rect -10850 15195 -10600 15255
rect -10850 15155 -10845 15195
rect -10805 15155 -10795 15195
rect -10755 15155 -10745 15195
rect -10705 15155 -10695 15195
rect -10655 15155 -10645 15195
rect -10605 15155 -10600 15195
rect -10850 15095 -10600 15155
rect -10850 15055 -10845 15095
rect -10805 15055 -10795 15095
rect -10755 15055 -10745 15095
rect -10705 15055 -10695 15095
rect -10655 15055 -10645 15095
rect -10605 15055 -10600 15095
rect -10850 14995 -10600 15055
rect -10850 14955 -10845 14995
rect -10805 14955 -10795 14995
rect -10755 14955 -10745 14995
rect -10705 14955 -10695 14995
rect -10655 14955 -10645 14995
rect -10605 14955 -10600 14995
rect -10850 14895 -10600 14955
rect -10850 14855 -10845 14895
rect -10805 14855 -10795 14895
rect -10755 14855 -10745 14895
rect -10705 14855 -10695 14895
rect -10655 14855 -10645 14895
rect -10605 14855 -10600 14895
rect -10850 14795 -10600 14855
rect -10850 14755 -10845 14795
rect -10805 14755 -10795 14795
rect -10755 14755 -10745 14795
rect -10705 14755 -10695 14795
rect -10655 14755 -10645 14795
rect -10605 14755 -10600 14795
rect -10850 14695 -10600 14755
rect -10850 14655 -10845 14695
rect -10805 14655 -10795 14695
rect -10755 14655 -10745 14695
rect -10705 14655 -10695 14695
rect -10655 14655 -10645 14695
rect -10605 14655 -10600 14695
rect -10850 12295 -10600 14655
rect -10850 12255 -10845 12295
rect -10805 12255 -10795 12295
rect -10755 12255 -10745 12295
rect -10705 12255 -10695 12295
rect -10655 12255 -10645 12295
rect -10605 12255 -10600 12295
rect -10850 12195 -10600 12255
rect -10850 12155 -10845 12195
rect -10805 12155 -10795 12195
rect -10755 12155 -10745 12195
rect -10705 12155 -10695 12195
rect -10655 12155 -10645 12195
rect -10605 12155 -10600 12195
rect -10850 12095 -10600 12155
rect -10850 12055 -10845 12095
rect -10805 12055 -10795 12095
rect -10755 12055 -10745 12095
rect -10705 12055 -10695 12095
rect -10655 12055 -10645 12095
rect -10605 12055 -10600 12095
rect -10850 11995 -10600 12055
rect -10850 11955 -10845 11995
rect -10805 11955 -10795 11995
rect -10755 11955 -10745 11995
rect -10705 11955 -10695 11995
rect -10655 11955 -10645 11995
rect -10605 11955 -10600 11995
rect -10850 11895 -10600 11955
rect -10850 11855 -10845 11895
rect -10805 11855 -10795 11895
rect -10755 11855 -10745 11895
rect -10705 11855 -10695 11895
rect -10655 11855 -10645 11895
rect -10605 11855 -10600 11895
rect -10850 11795 -10600 11855
rect -10850 11755 -10845 11795
rect -10805 11755 -10795 11795
rect -10755 11755 -10745 11795
rect -10705 11755 -10695 11795
rect -10655 11755 -10645 11795
rect -10605 11755 -10600 11795
rect -10850 11695 -10600 11755
rect -10850 11655 -10845 11695
rect -10805 11655 -10795 11695
rect -10755 11655 -10745 11695
rect -10705 11655 -10695 11695
rect -10655 11655 -10645 11695
rect -10605 11655 -10600 11695
rect -10850 11445 -10600 11655
rect -10850 11405 -10845 11445
rect -10805 11405 -10795 11445
rect -10755 11405 -10745 11445
rect -10705 11405 -10695 11445
rect -10655 11405 -10645 11445
rect -10605 11405 -10600 11445
rect -10850 11345 -10600 11405
rect -10850 11305 -10845 11345
rect -10805 11305 -10795 11345
rect -10755 11305 -10745 11345
rect -10705 11305 -10695 11345
rect -10655 11305 -10645 11345
rect -10605 11305 -10600 11345
rect -10850 11245 -10600 11305
rect -10850 11205 -10845 11245
rect -10805 11205 -10795 11245
rect -10755 11205 -10745 11245
rect -10705 11205 -10695 11245
rect -10655 11205 -10645 11245
rect -10605 11205 -10600 11245
rect -10850 11145 -10600 11205
rect -10850 11105 -10845 11145
rect -10805 11105 -10795 11145
rect -10755 11105 -10745 11145
rect -10705 11105 -10695 11145
rect -10655 11105 -10645 11145
rect -10605 11105 -10600 11145
rect -10850 11045 -10600 11105
rect -10850 11005 -10845 11045
rect -10805 11005 -10795 11045
rect -10755 11005 -10745 11045
rect -10705 11005 -10695 11045
rect -10655 11005 -10645 11045
rect -10605 11005 -10600 11045
rect -10850 10945 -10600 11005
rect -10850 10905 -10845 10945
rect -10805 10905 -10795 10945
rect -10755 10905 -10745 10945
rect -10705 10905 -10695 10945
rect -10655 10905 -10645 10945
rect -10605 10905 -10600 10945
rect -10850 10845 -10600 10905
rect -10850 10805 -10845 10845
rect -10805 10805 -10795 10845
rect -10755 10805 -10745 10845
rect -10705 10805 -10695 10845
rect -10655 10805 -10645 10845
rect -10605 10805 -10600 10845
rect -10850 8445 -10600 10805
rect -10850 8405 -10845 8445
rect -10805 8405 -10795 8445
rect -10755 8405 -10745 8445
rect -10705 8405 -10695 8445
rect -10655 8405 -10645 8445
rect -10605 8405 -10600 8445
rect -10850 8345 -10600 8405
rect -10850 8305 -10845 8345
rect -10805 8305 -10795 8345
rect -10755 8305 -10745 8345
rect -10705 8305 -10695 8345
rect -10655 8305 -10645 8345
rect -10605 8305 -10600 8345
rect -10850 8245 -10600 8305
rect -10850 8205 -10845 8245
rect -10805 8205 -10795 8245
rect -10755 8205 -10745 8245
rect -10705 8205 -10695 8245
rect -10655 8205 -10645 8245
rect -10605 8205 -10600 8245
rect -10850 8145 -10600 8205
rect -10850 8105 -10845 8145
rect -10805 8105 -10795 8145
rect -10755 8105 -10745 8145
rect -10705 8105 -10695 8145
rect -10655 8105 -10645 8145
rect -10605 8105 -10600 8145
rect -10850 8045 -10600 8105
rect -10850 8005 -10845 8045
rect -10805 8005 -10795 8045
rect -10755 8005 -10745 8045
rect -10705 8005 -10695 8045
rect -10655 8005 -10645 8045
rect -10605 8005 -10600 8045
rect -10850 7945 -10600 8005
rect -10850 7905 -10845 7945
rect -10805 7905 -10795 7945
rect -10755 7905 -10745 7945
rect -10705 7905 -10695 7945
rect -10655 7905 -10645 7945
rect -10605 7905 -10600 7945
rect -10850 7845 -10600 7905
rect -10850 7805 -10845 7845
rect -10805 7805 -10795 7845
rect -10755 7805 -10745 7845
rect -10705 7805 -10695 7845
rect -10655 7805 -10645 7845
rect -10605 7805 -10600 7845
rect -10850 7700 -10600 7805
rect -10550 14395 -10500 15400
rect -10550 14355 -10545 14395
rect -10505 14355 -10500 14395
rect -10550 13995 -10500 14355
rect -10550 13955 -10545 13995
rect -10505 13955 -10500 13995
rect -10550 13895 -10500 13955
rect -10550 13855 -10545 13895
rect -10505 13855 -10500 13895
rect -10550 13795 -10500 13855
rect -10550 13755 -10545 13795
rect -10505 13755 -10500 13795
rect -10550 13595 -10500 13755
rect -10550 13555 -10545 13595
rect -10505 13555 -10500 13595
rect -10550 13395 -10500 13555
rect -10550 13355 -10545 13395
rect -10505 13355 -10500 13395
rect -10550 13195 -10500 13355
rect -10550 13155 -10545 13195
rect -10505 13155 -10500 13195
rect -10550 13095 -10500 13155
rect -10550 13055 -10545 13095
rect -10505 13055 -10500 13095
rect -10550 12995 -10500 13055
rect -10550 12955 -10545 12995
rect -10505 12955 -10500 12995
rect -10550 12595 -10500 12955
rect -10550 12555 -10545 12595
rect -10505 12555 -10500 12595
rect -10550 10545 -10500 12555
rect -10550 10505 -10545 10545
rect -10505 10505 -10500 10545
rect -10550 10145 -10500 10505
rect -10550 10105 -10545 10145
rect -10505 10105 -10500 10145
rect -10550 10045 -10500 10105
rect -10550 10005 -10545 10045
rect -10505 10005 -10500 10045
rect -10550 9945 -10500 10005
rect -10550 9905 -10545 9945
rect -10505 9905 -10500 9945
rect -10550 9745 -10500 9905
rect -10550 9705 -10545 9745
rect -10505 9705 -10500 9745
rect -10550 9545 -10500 9705
rect -10550 9505 -10545 9545
rect -10505 9505 -10500 9545
rect -10550 9345 -10500 9505
rect -10550 9305 -10545 9345
rect -10505 9305 -10500 9345
rect -10550 9245 -10500 9305
rect -10550 9205 -10545 9245
rect -10505 9205 -10500 9245
rect -10550 9145 -10500 9205
rect -10550 9105 -10545 9145
rect -10505 9105 -10500 9145
rect -10550 8745 -10500 9105
rect -10550 8705 -10545 8745
rect -10505 8705 -10500 8745
rect -10550 7700 -10500 8705
rect -10450 13295 -10400 15400
rect -10450 13255 -10445 13295
rect -10405 13255 -10400 13295
rect -10450 7700 -10400 13255
rect -10350 14395 -10300 15400
rect -10350 14355 -10345 14395
rect -10305 14355 -10300 14395
rect -10350 13995 -10300 14355
rect -10350 13955 -10345 13995
rect -10305 13955 -10300 13995
rect -10350 13895 -10300 13955
rect -10350 13855 -10345 13895
rect -10305 13855 -10300 13895
rect -10350 13795 -10300 13855
rect -10350 13755 -10345 13795
rect -10305 13755 -10300 13795
rect -10350 13595 -10300 13755
rect -10350 13555 -10345 13595
rect -10305 13555 -10300 13595
rect -10350 13395 -10300 13555
rect -10350 13355 -10345 13395
rect -10305 13355 -10300 13395
rect -10350 13195 -10300 13355
rect -10350 13155 -10345 13195
rect -10305 13155 -10300 13195
rect -10350 13095 -10300 13155
rect -10350 13055 -10345 13095
rect -10305 13055 -10300 13095
rect -10350 12995 -10300 13055
rect -10350 12955 -10345 12995
rect -10305 12955 -10300 12995
rect -10350 12595 -10300 12955
rect -10350 12555 -10345 12595
rect -10305 12555 -10300 12595
rect -10350 10545 -10300 12555
rect -10350 10505 -10345 10545
rect -10305 10505 -10300 10545
rect -10350 10145 -10300 10505
rect -10350 10105 -10345 10145
rect -10305 10105 -10300 10145
rect -10350 10045 -10300 10105
rect -10350 10005 -10345 10045
rect -10305 10005 -10300 10045
rect -10350 9945 -10300 10005
rect -10350 9905 -10345 9945
rect -10305 9905 -10300 9945
rect -10350 9745 -10300 9905
rect -10350 9705 -10345 9745
rect -10305 9705 -10300 9745
rect -10350 9545 -10300 9705
rect -10350 9505 -10345 9545
rect -10305 9505 -10300 9545
rect -10350 9345 -10300 9505
rect -10350 9305 -10345 9345
rect -10305 9305 -10300 9345
rect -10350 9245 -10300 9305
rect -10350 9205 -10345 9245
rect -10305 9205 -10300 9245
rect -10350 9145 -10300 9205
rect -10350 9105 -10345 9145
rect -10305 9105 -10300 9145
rect -10350 8745 -10300 9105
rect -10350 8705 -10345 8745
rect -10305 8705 -10300 8745
rect -10350 7700 -10300 8705
rect -10250 13695 -10200 15400
rect -10250 13655 -10245 13695
rect -10205 13655 -10200 13695
rect -10250 7700 -10200 13655
rect -10150 14395 -10100 15400
rect -10150 14355 -10145 14395
rect -10105 14355 -10100 14395
rect -10150 13995 -10100 14355
rect -10150 13955 -10145 13995
rect -10105 13955 -10100 13995
rect -10150 13895 -10100 13955
rect -10150 13855 -10145 13895
rect -10105 13855 -10100 13895
rect -10150 13795 -10100 13855
rect -10150 13755 -10145 13795
rect -10105 13755 -10100 13795
rect -10150 13595 -10100 13755
rect -10150 13555 -10145 13595
rect -10105 13555 -10100 13595
rect -10150 13395 -10100 13555
rect -10150 13355 -10145 13395
rect -10105 13355 -10100 13395
rect -10150 13195 -10100 13355
rect -10150 13155 -10145 13195
rect -10105 13155 -10100 13195
rect -10150 13095 -10100 13155
rect -10150 13055 -10145 13095
rect -10105 13055 -10100 13095
rect -10150 12995 -10100 13055
rect -10150 12955 -10145 12995
rect -10105 12955 -10100 12995
rect -10150 12595 -10100 12955
rect -10150 12555 -10145 12595
rect -10105 12555 -10100 12595
rect -10150 10545 -10100 12555
rect -10150 10505 -10145 10545
rect -10105 10505 -10100 10545
rect -10150 10145 -10100 10505
rect -10150 10105 -10145 10145
rect -10105 10105 -10100 10145
rect -10150 10045 -10100 10105
rect -10150 10005 -10145 10045
rect -10105 10005 -10100 10045
rect -10150 9945 -10100 10005
rect -10150 9905 -10145 9945
rect -10105 9905 -10100 9945
rect -10150 9745 -10100 9905
rect -10150 9705 -10145 9745
rect -10105 9705 -10100 9745
rect -10150 9545 -10100 9705
rect -10150 9505 -10145 9545
rect -10105 9505 -10100 9545
rect -10150 9345 -10100 9505
rect -10150 9305 -10145 9345
rect -10105 9305 -10100 9345
rect -10150 9245 -10100 9305
rect -10150 9205 -10145 9245
rect -10105 9205 -10100 9245
rect -10150 9145 -10100 9205
rect -10150 9105 -10145 9145
rect -10105 9105 -10100 9145
rect -10150 8745 -10100 9105
rect -10150 8705 -10145 8745
rect -10105 8705 -10100 8745
rect -10150 7700 -10100 8705
rect -10050 9845 -10000 15400
rect -10050 9805 -10045 9845
rect -10005 9805 -10000 9845
rect -10050 7700 -10000 9805
rect -9950 14395 -9900 15400
rect -9950 14355 -9945 14395
rect -9905 14355 -9900 14395
rect -9950 13995 -9900 14355
rect -9950 13955 -9945 13995
rect -9905 13955 -9900 13995
rect -9950 13895 -9900 13955
rect -9950 13855 -9945 13895
rect -9905 13855 -9900 13895
rect -9950 13795 -9900 13855
rect -9950 13755 -9945 13795
rect -9905 13755 -9900 13795
rect -9950 13595 -9900 13755
rect -9950 13555 -9945 13595
rect -9905 13555 -9900 13595
rect -9950 13395 -9900 13555
rect -9950 13355 -9945 13395
rect -9905 13355 -9900 13395
rect -9950 13195 -9900 13355
rect -9950 13155 -9945 13195
rect -9905 13155 -9900 13195
rect -9950 13095 -9900 13155
rect -9950 13055 -9945 13095
rect -9905 13055 -9900 13095
rect -9950 12995 -9900 13055
rect -9950 12955 -9945 12995
rect -9905 12955 -9900 12995
rect -9950 12595 -9900 12955
rect -9950 12555 -9945 12595
rect -9905 12555 -9900 12595
rect -9950 10545 -9900 12555
rect -9950 10505 -9945 10545
rect -9905 10505 -9900 10545
rect -9950 10145 -9900 10505
rect -9950 10105 -9945 10145
rect -9905 10105 -9900 10145
rect -9950 10045 -9900 10105
rect -9950 10005 -9945 10045
rect -9905 10005 -9900 10045
rect -9950 9945 -9900 10005
rect -9950 9905 -9945 9945
rect -9905 9905 -9900 9945
rect -9950 9745 -9900 9905
rect -9950 9705 -9945 9745
rect -9905 9705 -9900 9745
rect -9950 9545 -9900 9705
rect -9950 9505 -9945 9545
rect -9905 9505 -9900 9545
rect -9950 9345 -9900 9505
rect -9950 9305 -9945 9345
rect -9905 9305 -9900 9345
rect -9950 9245 -9900 9305
rect -9950 9205 -9945 9245
rect -9905 9205 -9900 9245
rect -9950 9145 -9900 9205
rect -9950 9105 -9945 9145
rect -9905 9105 -9900 9145
rect -9950 8745 -9900 9105
rect -9950 8705 -9945 8745
rect -9905 8705 -9900 8745
rect -9950 7700 -9900 8705
rect -9850 9445 -9800 15400
rect -9850 9405 -9845 9445
rect -9805 9405 -9800 9445
rect -9850 7700 -9800 9405
rect -9750 14395 -9700 15400
rect -9750 14355 -9745 14395
rect -9705 14355 -9700 14395
rect -9750 13995 -9700 14355
rect -9750 13955 -9745 13995
rect -9705 13955 -9700 13995
rect -9750 13895 -9700 13955
rect -9750 13855 -9745 13895
rect -9705 13855 -9700 13895
rect -9750 13795 -9700 13855
rect -9750 13755 -9745 13795
rect -9705 13755 -9700 13795
rect -9750 13595 -9700 13755
rect -9750 13555 -9745 13595
rect -9705 13555 -9700 13595
rect -9750 13395 -9700 13555
rect -9750 13355 -9745 13395
rect -9705 13355 -9700 13395
rect -9750 13195 -9700 13355
rect -9750 13155 -9745 13195
rect -9705 13155 -9700 13195
rect -9750 13095 -9700 13155
rect -9750 13055 -9745 13095
rect -9705 13055 -9700 13095
rect -9750 12995 -9700 13055
rect -9750 12955 -9745 12995
rect -9705 12955 -9700 12995
rect -9750 12595 -9700 12955
rect -9750 12555 -9745 12595
rect -9705 12555 -9700 12595
rect -9750 10545 -9700 12555
rect -9750 10505 -9745 10545
rect -9705 10505 -9700 10545
rect -9750 10145 -9700 10505
rect -9750 10105 -9745 10145
rect -9705 10105 -9700 10145
rect -9750 10045 -9700 10105
rect -9750 10005 -9745 10045
rect -9705 10005 -9700 10045
rect -9750 9945 -9700 10005
rect -9750 9905 -9745 9945
rect -9705 9905 -9700 9945
rect -9750 9745 -9700 9905
rect -9750 9705 -9745 9745
rect -9705 9705 -9700 9745
rect -9750 9545 -9700 9705
rect -9750 9505 -9745 9545
rect -9705 9505 -9700 9545
rect -9750 9345 -9700 9505
rect -9750 9305 -9745 9345
rect -9705 9305 -9700 9345
rect -9750 9245 -9700 9305
rect -9750 9205 -9745 9245
rect -9705 9205 -9700 9245
rect -9750 9145 -9700 9205
rect -9750 9105 -9745 9145
rect -9705 9105 -9700 9145
rect -9750 8745 -9700 9105
rect -9750 8705 -9745 8745
rect -9705 8705 -9700 8745
rect -9750 7700 -9700 8705
rect -9500 13495 -9450 15400
rect -9500 13455 -9495 13495
rect -9455 13455 -9450 13495
rect -9500 9645 -9450 13455
rect -9500 9605 -9495 9645
rect -9455 9605 -9450 9645
rect -9500 7700 -9450 9605
rect -9350 13495 -9300 15400
rect -9350 13455 -9345 13495
rect -9305 13455 -9300 13495
rect -9350 9645 -9300 13455
rect -9350 9605 -9345 9645
rect -9305 9605 -9300 9645
rect -9350 7700 -9300 9605
rect 13250 14395 13300 15400
rect 13250 14355 13255 14395
rect 13295 14355 13300 14395
rect 13250 13995 13300 14355
rect 13250 13955 13255 13995
rect 13295 13955 13300 13995
rect 13250 13895 13300 13955
rect 13250 13855 13255 13895
rect 13295 13855 13300 13895
rect 13250 13795 13300 13855
rect 13250 13755 13255 13795
rect 13295 13755 13300 13795
rect 13250 13695 13300 13755
rect 13250 13655 13255 13695
rect 13295 13655 13300 13695
rect 13250 13595 13300 13655
rect 13250 13555 13255 13595
rect 13295 13555 13300 13595
rect 13250 13395 13300 13555
rect 13250 13355 13255 13395
rect 13295 13355 13300 13395
rect 13250 13295 13300 13355
rect 13250 13255 13255 13295
rect 13295 13255 13300 13295
rect 13250 13195 13300 13255
rect 13250 13155 13255 13195
rect 13295 13155 13300 13195
rect 13250 13095 13300 13155
rect 13250 13055 13255 13095
rect 13295 13055 13300 13095
rect 13250 12995 13300 13055
rect 13250 12955 13255 12995
rect 13295 12955 13300 12995
rect 13250 12595 13300 12955
rect 13250 12555 13255 12595
rect 13295 12555 13300 12595
rect 13250 11595 13300 12555
rect 13250 11555 13255 11595
rect 13295 11555 13300 11595
rect 13250 11545 13300 11555
rect 13250 11505 13255 11545
rect 13295 11505 13300 11545
rect 13250 10545 13300 11505
rect 13250 10505 13255 10545
rect 13295 10505 13300 10545
rect 13250 10145 13300 10505
rect 13250 10105 13255 10145
rect 13295 10105 13300 10145
rect 13250 10045 13300 10105
rect 13250 10005 13255 10045
rect 13295 10005 13300 10045
rect 13250 9945 13300 10005
rect 13250 9905 13255 9945
rect 13295 9905 13300 9945
rect 13250 9845 13300 9905
rect 13250 9805 13255 9845
rect 13295 9805 13300 9845
rect 13250 9745 13300 9805
rect 13250 9705 13255 9745
rect 13295 9705 13300 9745
rect 13250 9545 13300 9705
rect 13250 9505 13255 9545
rect 13295 9505 13300 9545
rect 13250 9445 13300 9505
rect 13250 9405 13255 9445
rect 13295 9405 13300 9445
rect 13250 9345 13300 9405
rect 13250 9305 13255 9345
rect 13295 9305 13300 9345
rect 13250 9245 13300 9305
rect 13250 9205 13255 9245
rect 13295 9205 13300 9245
rect 13250 9145 13300 9205
rect 13250 9105 13255 9145
rect 13295 9105 13300 9145
rect 13250 8745 13300 9105
rect 13250 8705 13255 8745
rect 13295 8705 13300 8745
rect 13250 7745 13300 8705
rect 13250 7705 13255 7745
rect 13295 7705 13300 7745
rect 13250 7700 13300 7705
rect 13350 14295 13400 15400
rect 13350 14255 13355 14295
rect 13395 14255 13400 14295
rect 13350 14095 13400 14255
rect 13350 14055 13355 14095
rect 13395 14055 13400 14095
rect 13350 11695 13400 14055
rect 13350 11655 13355 11695
rect 13395 11655 13400 11695
rect 13350 9045 13400 11655
rect 13350 9005 13355 9045
rect 13395 9005 13400 9045
rect 13350 8845 13400 9005
rect 13350 8805 13355 8845
rect 13395 8805 13400 8845
rect 13350 7700 13400 8805
rect 13450 14195 13500 15400
rect 13450 14155 13455 14195
rect 13495 14155 13500 14195
rect 13450 11895 13500 14155
rect 13450 11855 13455 11895
rect 13495 11855 13500 11895
rect 13450 8945 13500 11855
rect 13450 8905 13455 8945
rect 13495 8905 13500 8945
rect 13450 7700 13500 8905
rect 13550 14295 13600 15400
rect 13550 14255 13555 14295
rect 13595 14255 13600 14295
rect 13550 14095 13600 14255
rect 13550 14055 13555 14095
rect 13595 14055 13600 14095
rect 13550 11695 13600 14055
rect 13550 11655 13555 11695
rect 13595 11655 13600 11695
rect 13550 9045 13600 11655
rect 13550 9005 13555 9045
rect 13595 9005 13600 9045
rect 13550 8845 13600 9005
rect 13550 8805 13555 8845
rect 13595 8805 13600 8845
rect 13550 7700 13600 8805
rect 13650 14395 13700 15400
rect 13650 14355 13655 14395
rect 13695 14355 13700 14395
rect 13650 13995 13700 14355
rect 13650 13955 13655 13995
rect 13695 13955 13700 13995
rect 13650 13895 13700 13955
rect 13650 13855 13655 13895
rect 13695 13855 13700 13895
rect 13650 13795 13700 13855
rect 13650 13755 13655 13795
rect 13695 13755 13700 13795
rect 13650 13695 13700 13755
rect 13650 13655 13655 13695
rect 13695 13655 13700 13695
rect 13650 13595 13700 13655
rect 13650 13555 13655 13595
rect 13695 13555 13700 13595
rect 13650 13395 13700 13555
rect 13650 13355 13655 13395
rect 13695 13355 13700 13395
rect 13650 13295 13700 13355
rect 13650 13255 13655 13295
rect 13695 13255 13700 13295
rect 13650 13195 13700 13255
rect 13650 13155 13655 13195
rect 13695 13155 13700 13195
rect 13650 13095 13700 13155
rect 13650 13055 13655 13095
rect 13695 13055 13700 13095
rect 13650 12995 13700 13055
rect 13650 12955 13655 12995
rect 13695 12955 13700 12995
rect 13650 12595 13700 12955
rect 13650 12555 13655 12595
rect 13695 12555 13700 12595
rect 13650 11595 13700 12555
rect 13650 11555 13655 11595
rect 13695 11555 13700 11595
rect 13650 11545 13700 11555
rect 13650 11505 13655 11545
rect 13695 11505 13700 11545
rect 13650 10545 13700 11505
rect 13650 10505 13655 10545
rect 13695 10505 13700 10545
rect 13650 10145 13700 10505
rect 13650 10105 13655 10145
rect 13695 10105 13700 10145
rect 13650 10045 13700 10105
rect 13650 10005 13655 10045
rect 13695 10005 13700 10045
rect 13650 9945 13700 10005
rect 13650 9905 13655 9945
rect 13695 9905 13700 9945
rect 13650 9845 13700 9905
rect 13650 9805 13655 9845
rect 13695 9805 13700 9845
rect 13650 9745 13700 9805
rect 13650 9705 13655 9745
rect 13695 9705 13700 9745
rect 13650 9545 13700 9705
rect 13650 9505 13655 9545
rect 13695 9505 13700 9545
rect 13650 9445 13700 9505
rect 13650 9405 13655 9445
rect 13695 9405 13700 9445
rect 13650 9345 13700 9405
rect 13650 9305 13655 9345
rect 13695 9305 13700 9345
rect 13650 9245 13700 9305
rect 13650 9205 13655 9245
rect 13695 9205 13700 9245
rect 13650 9145 13700 9205
rect 13650 9105 13655 9145
rect 13695 9105 13700 9145
rect 13650 8745 13700 9105
rect 13650 8705 13655 8745
rect 13695 8705 13700 8745
rect 13650 7745 13700 8705
rect 13650 7705 13655 7745
rect 13695 7705 13700 7745
rect 13650 7700 13700 7705
rect 13750 12895 13800 15400
rect 13750 12855 13755 12895
rect 13795 12855 13800 12895
rect 13750 12695 13800 12855
rect 13750 12655 13755 12695
rect 13795 12655 13800 12695
rect 13750 11445 13800 12655
rect 13750 11405 13755 11445
rect 13795 11405 13800 11445
rect 13750 10445 13800 11405
rect 13750 10405 13755 10445
rect 13795 10405 13800 10445
rect 13750 10245 13800 10405
rect 13750 10205 13755 10245
rect 13795 10205 13800 10245
rect 13750 7700 13800 10205
rect 13850 12795 13900 15400
rect 13850 12755 13855 12795
rect 13895 12755 13900 12795
rect 13850 11245 13900 12755
rect 13850 11205 13855 11245
rect 13895 11205 13900 11245
rect 13850 10345 13900 11205
rect 13850 10305 13855 10345
rect 13895 10305 13900 10345
rect 13850 7700 13900 10305
rect 13950 12895 14000 15400
rect 13950 12855 13955 12895
rect 13995 12855 14000 12895
rect 13950 12695 14000 12855
rect 13950 12655 13955 12695
rect 13995 12655 14000 12695
rect 13950 11445 14000 12655
rect 14050 15395 14100 15400
rect 14050 15355 14055 15395
rect 14095 15355 14100 15395
rect 14050 11950 14100 15355
rect 21900 15395 21950 15400
rect 21900 15355 21905 15395
rect 21945 15355 21950 15395
rect 14150 15200 21850 15300
rect 14150 11950 14250 15200
rect 21750 11950 21850 15200
rect 14150 11900 21850 11950
rect 14050 11895 21850 11900
rect 14050 11855 14055 11895
rect 14095 11855 21850 11895
rect 14050 11850 21850 11855
rect 13950 11405 13955 11445
rect 13995 11405 14000 11445
rect 13950 10445 14000 11405
rect 14050 11595 14100 11800
rect 14150 11795 21850 11800
rect 14150 11755 14155 11795
rect 14195 11755 14205 11795
rect 14245 11755 14255 11795
rect 14295 11755 14305 11795
rect 14345 11755 14355 11795
rect 14395 11755 14405 11795
rect 14445 11755 14455 11795
rect 14495 11755 14505 11795
rect 14545 11755 14555 11795
rect 14595 11755 14605 11795
rect 14645 11755 14655 11795
rect 14695 11755 14705 11795
rect 14745 11755 14755 11795
rect 14795 11755 14805 11795
rect 14845 11755 14855 11795
rect 14895 11755 14905 11795
rect 14945 11755 14955 11795
rect 14995 11755 15005 11795
rect 15045 11755 15055 11795
rect 15095 11755 15105 11795
rect 15145 11755 15155 11795
rect 15195 11755 15205 11795
rect 15245 11755 15255 11795
rect 15295 11755 15305 11795
rect 15345 11755 15355 11795
rect 15395 11755 15405 11795
rect 15445 11755 15455 11795
rect 15495 11755 15505 11795
rect 15545 11755 15555 11795
rect 15595 11755 15605 11795
rect 15645 11755 15655 11795
rect 15695 11755 15705 11795
rect 15745 11755 15755 11795
rect 15795 11755 15805 11795
rect 15845 11755 15855 11795
rect 15895 11755 15905 11795
rect 15945 11755 15955 11795
rect 15995 11755 16005 11795
rect 16045 11755 16055 11795
rect 16095 11755 16105 11795
rect 16145 11755 16155 11795
rect 16195 11755 16205 11795
rect 16245 11755 16255 11795
rect 16295 11755 16305 11795
rect 16345 11755 16355 11795
rect 16395 11755 16405 11795
rect 16445 11755 16455 11795
rect 16495 11755 16505 11795
rect 16545 11755 16555 11795
rect 16595 11755 16605 11795
rect 16645 11755 16655 11795
rect 16695 11755 21705 11795
rect 21745 11755 21755 11795
rect 21795 11755 21805 11795
rect 21845 11755 21850 11795
rect 14150 11695 21850 11755
rect 14150 11655 14155 11695
rect 14195 11655 14205 11695
rect 14245 11655 14255 11695
rect 14295 11655 14305 11695
rect 14345 11655 14355 11695
rect 14395 11655 14405 11695
rect 14445 11655 14455 11695
rect 14495 11655 14505 11695
rect 14545 11655 14555 11695
rect 14595 11655 14605 11695
rect 14645 11655 14655 11695
rect 14695 11655 14705 11695
rect 14745 11655 14755 11695
rect 14795 11655 14805 11695
rect 14845 11655 14855 11695
rect 14895 11655 14905 11695
rect 14945 11655 14955 11695
rect 14995 11655 15005 11695
rect 15045 11655 15055 11695
rect 15095 11655 15105 11695
rect 15145 11655 15155 11695
rect 15195 11655 15205 11695
rect 15245 11655 15255 11695
rect 15295 11655 15305 11695
rect 15345 11655 15355 11695
rect 15395 11655 15405 11695
rect 15445 11655 15455 11695
rect 15495 11655 15505 11695
rect 15545 11655 15555 11695
rect 15595 11655 15605 11695
rect 15645 11655 15655 11695
rect 15695 11655 15705 11695
rect 15745 11655 15755 11695
rect 15795 11655 15805 11695
rect 15845 11655 15855 11695
rect 15895 11655 15905 11695
rect 15945 11655 15955 11695
rect 15995 11655 16005 11695
rect 16045 11655 16055 11695
rect 16095 11655 16105 11695
rect 16145 11655 16155 11695
rect 16195 11655 16205 11695
rect 16245 11655 16255 11695
rect 16295 11655 16305 11695
rect 16345 11655 16355 11695
rect 16395 11655 16405 11695
rect 16445 11655 16455 11695
rect 16495 11655 16505 11695
rect 16545 11655 16555 11695
rect 16595 11655 16605 11695
rect 16645 11655 16655 11695
rect 16695 11655 21705 11695
rect 21745 11655 21755 11695
rect 21795 11655 21805 11695
rect 21845 11655 21850 11695
rect 14150 11650 21850 11655
rect 14050 11555 14055 11595
rect 14095 11555 14100 11595
rect 14050 11545 14100 11555
rect 14050 11505 14055 11545
rect 14095 11505 14100 11545
rect 14050 11300 14100 11505
rect 21900 11595 21950 15355
rect 21900 11555 21905 11595
rect 21945 11555 21950 11595
rect 21900 11545 21950 11555
rect 21900 11505 21905 11545
rect 21945 11505 21950 11545
rect 14150 11445 21850 11450
rect 14150 11405 14155 11445
rect 14195 11405 14205 11445
rect 14245 11405 14255 11445
rect 14295 11405 14305 11445
rect 14345 11405 14355 11445
rect 14395 11405 14405 11445
rect 14445 11405 14455 11445
rect 14495 11405 14505 11445
rect 14545 11405 14555 11445
rect 14595 11405 14605 11445
rect 14645 11405 14655 11445
rect 14695 11405 14705 11445
rect 14745 11405 14755 11445
rect 14795 11405 14805 11445
rect 14845 11405 14855 11445
rect 14895 11405 14905 11445
rect 14945 11405 14955 11445
rect 14995 11405 15005 11445
rect 15045 11405 15055 11445
rect 15095 11405 15105 11445
rect 15145 11405 15155 11445
rect 15195 11405 15205 11445
rect 15245 11405 15255 11445
rect 15295 11405 15305 11445
rect 15345 11405 15355 11445
rect 15395 11405 15405 11445
rect 15445 11405 15455 11445
rect 15495 11405 15505 11445
rect 15545 11405 15555 11445
rect 15595 11405 15605 11445
rect 15645 11405 15655 11445
rect 15695 11405 15705 11445
rect 15745 11405 15755 11445
rect 15795 11405 15805 11445
rect 15845 11405 15855 11445
rect 15895 11405 15905 11445
rect 15945 11405 15955 11445
rect 15995 11405 16005 11445
rect 16045 11405 16055 11445
rect 16095 11405 16105 11445
rect 16145 11405 16155 11445
rect 16195 11405 16205 11445
rect 16245 11405 16255 11445
rect 16295 11405 16305 11445
rect 16345 11405 16355 11445
rect 16395 11405 16405 11445
rect 16445 11405 16455 11445
rect 16495 11405 16505 11445
rect 16545 11405 16555 11445
rect 16595 11405 16605 11445
rect 16645 11405 16655 11445
rect 16695 11405 21705 11445
rect 21745 11405 21755 11445
rect 21795 11405 21805 11445
rect 21845 11405 21850 11445
rect 14150 11345 21850 11405
rect 14150 11305 14155 11345
rect 14195 11305 14205 11345
rect 14245 11305 14255 11345
rect 14295 11305 14305 11345
rect 14345 11305 14355 11345
rect 14395 11305 14405 11345
rect 14445 11305 14455 11345
rect 14495 11305 14505 11345
rect 14545 11305 14555 11345
rect 14595 11305 14605 11345
rect 14645 11305 14655 11345
rect 14695 11305 14705 11345
rect 14745 11305 14755 11345
rect 14795 11305 14805 11345
rect 14845 11305 14855 11345
rect 14895 11305 14905 11345
rect 14945 11305 14955 11345
rect 14995 11305 15005 11345
rect 15045 11305 15055 11345
rect 15095 11305 15105 11345
rect 15145 11305 15155 11345
rect 15195 11305 15205 11345
rect 15245 11305 15255 11345
rect 15295 11305 15305 11345
rect 15345 11305 15355 11345
rect 15395 11305 15405 11345
rect 15445 11305 15455 11345
rect 15495 11305 15505 11345
rect 15545 11305 15555 11345
rect 15595 11305 15605 11345
rect 15645 11305 15655 11345
rect 15695 11305 15705 11345
rect 15745 11305 15755 11345
rect 15795 11305 15805 11345
rect 15845 11305 15855 11345
rect 15895 11305 15905 11345
rect 15945 11305 15955 11345
rect 15995 11305 16005 11345
rect 16045 11305 16055 11345
rect 16095 11305 16105 11345
rect 16145 11305 16155 11345
rect 16195 11305 16205 11345
rect 16245 11305 16255 11345
rect 16295 11305 16305 11345
rect 16345 11305 16355 11345
rect 16395 11305 16405 11345
rect 16445 11305 16455 11345
rect 16495 11305 16505 11345
rect 16545 11305 16555 11345
rect 16595 11305 16605 11345
rect 16645 11305 16655 11345
rect 16695 11305 21705 11345
rect 21745 11305 21755 11345
rect 21795 11305 21805 11345
rect 21845 11305 21850 11345
rect 14150 11300 21850 11305
rect 14050 11245 21850 11250
rect 14050 11205 14055 11245
rect 14095 11205 21850 11245
rect 14050 11200 21850 11205
rect 14150 11150 21850 11200
rect 13950 10405 13955 10445
rect 13995 10405 14000 10445
rect 13950 10245 14000 10405
rect 13950 10205 13955 10245
rect 13995 10205 14000 10245
rect 13950 7700 14000 10205
rect 14050 8745 14100 11150
rect 14050 8705 14055 8745
rect 14095 8705 14100 8745
rect 14050 7700 14100 8705
rect 14150 7900 14250 11150
rect 21750 7900 21850 11150
rect 14150 7800 21850 7900
rect 21900 7745 21950 11505
rect 21900 7705 21905 7745
rect 21945 7705 21950 7745
rect 21900 7700 21950 7705
use ddab_slice  ddab_slice_0
timestamp 1726832924
transform -1 0 5450 0 -1 15400
box -7200 0 14550 7700
use invdummy  invdummy_0
timestamp 1722856725
transform 1 0 12550 0 1 11550
box -50 0 300 3850
use invdummy  invdummy_3
timestamp 1722856725
transform 1 0 12550 0 1 7700
box -50 0 300 3850
use invdummy  invdummy_5
timestamp 1722856725
transform -1 0 -9000 0 1 11550
box -50 0 300 3850
use invdummy  invdummy_7
timestamp 1722856725
transform -1 0 -9000 0 1 7700
box -50 0 300 3850
use invedge  invedge_0
timestamp 1722865417
transform 1 0 12600 0 1 10450
box 150 1100 600 4950
use invedge  invedge_3
timestamp 1722865417
transform 1 0 12600 0 1 6600
box 150 1100 600 4950
use invedge  invedge_5
timestamp 1722865417
transform -1 0 -9050 0 1 10450
box 150 1100 600 4950
use invedge  invedge_7
timestamp 1722865417
transform -1 0 -9050 0 1 6600
box 150 1100 600 4950
<< labels >>
rlabel metal4 -10450 15350 -10400 15400 0 ipa
port 1 nsew
rlabel metal4 -10250 15350 -10200 15400 0 ima
port 2 nsew
rlabel metal4 -10050 15350 -10000 15400 0 ipb
port 3 nsew
rlabel metal4 -9850 15350 -9800 15400 0 imb
port 4 nsew
rlabel metal4 -9500 15350 -9450 15400 0 bp
port 7 nsew
rlabel metal4 -9350 15350 -9300 15400 0 bn
port 8 nsew
rlabel metal4 -10850 15350 -10600 15400 0 vdd
port 9 nsew
rlabel metal4 -10550 15350 -10500 15400 0 vss
port 10 nsew
rlabel metal4 -10950 15350 -10900 15400 0 vsub
port 11 nsew
rlabel metal4 13750 15350 13800 15400 0 op
port 5 nsew
rlabel metal4 13950 15350 14000 15400 0 op
port 5 nsew
rlabel metal4 13350 15350 13400 15400 0 om
port 6 nsew
rlabel metal4 13550 15350 13600 15400 0 om
port 6 nsew
rlabel metal4 13850 15350 13900 15400 0 xm
rlabel metal4 13450 15350 13500 15400 0 xp
<< end >>
