magic
tech sky130A
timestamp 1726842748
<< locali >>
rect 150 13485 200 13500
rect 150 13465 165 13485
rect 185 13465 200 13485
rect 150 13450 200 13465
rect 300 13485 350 13500
rect 300 13465 315 13485
rect 335 13465 350 13485
rect 300 13450 350 13465
rect 150 9635 200 9650
rect 150 9615 165 9635
rect 185 9615 200 9635
rect 150 9600 200 9615
rect 300 9635 350 9650
rect 300 9615 315 9635
rect 335 9615 350 9635
rect 300 9600 350 9615
<< viali >>
rect 165 13465 185 13485
rect 315 13465 335 13485
rect 15 11565 35 11585
rect 15 11515 35 11535
rect 165 9615 185 9635
rect 315 9615 335 9635
<< metal1 >>
rect 150 13490 200 13500
rect 150 13460 160 13490
rect 190 13460 200 13490
rect 150 13450 200 13460
rect 300 13490 350 13500
rect 300 13460 310 13490
rect 340 13460 350 13490
rect 300 13450 350 13460
rect 0 11590 50 11600
rect 0 11560 10 11590
rect 40 11560 50 11590
rect 0 11540 50 11560
rect 0 11510 10 11540
rect 40 11510 50 11540
rect 0 11500 50 11510
rect 150 9640 200 9650
rect 150 9610 160 9640
rect 190 9610 200 9640
rect 150 9600 200 9610
rect 300 9640 350 9650
rect 300 9610 310 9640
rect 340 9610 350 9640
rect 300 9600 350 9610
<< via1 >>
rect 160 13485 190 13490
rect 160 13465 165 13485
rect 165 13465 185 13485
rect 185 13465 190 13485
rect 160 13460 190 13465
rect 310 13485 340 13490
rect 310 13465 315 13485
rect 315 13465 335 13485
rect 335 13465 340 13485
rect 310 13460 340 13465
rect 10 11585 40 11590
rect 10 11565 15 11585
rect 15 11565 35 11585
rect 35 11565 40 11585
rect 10 11560 40 11565
rect 10 11535 40 11540
rect 10 11515 15 11535
rect 15 11515 35 11535
rect 35 11515 40 11535
rect 10 11510 40 11515
rect 160 9635 190 9640
rect 160 9615 165 9635
rect 165 9615 185 9635
rect 185 9615 190 9635
rect 160 9610 190 9615
rect 310 9635 340 9640
rect 310 9615 315 9635
rect 315 9615 335 9635
rect 335 9615 340 9635
rect 310 9610 340 9615
<< metal2 >>
rect 150 13490 200 13500
rect 150 13460 160 13490
rect 190 13460 200 13490
rect 150 13450 200 13460
rect 300 13490 350 13500
rect 300 13460 310 13490
rect 340 13460 350 13490
rect 300 13450 350 13460
rect 0 11590 50 11600
rect 0 11560 10 11590
rect 40 11560 50 11590
rect 0 11540 50 11560
rect 0 11510 10 11540
rect 40 11510 50 11540
rect 0 11500 50 11510
rect 150 9640 200 9650
rect 150 9610 160 9640
rect 190 9610 200 9640
rect 150 9600 200 9610
rect 300 9640 350 9650
rect 300 9610 310 9640
rect 340 9610 350 9640
rect 300 9600 350 9610
<< via2 >>
rect 160 13460 190 13490
rect 310 13460 340 13490
rect 10 11560 40 11590
rect 10 11510 40 11540
rect 160 9610 190 9640
rect 310 9610 340 9640
<< metal3 >>
rect -1200 15295 0 15300
rect -1200 15255 -1195 15295
rect -1155 15255 -1145 15295
rect -1105 15255 -1095 15295
rect -1055 15255 -1045 15295
rect -1005 15255 -995 15295
rect -955 15255 0 15295
rect -1200 15250 0 15255
rect 22850 15295 24050 15300
rect 22850 15255 23805 15295
rect 23845 15255 23855 15295
rect 23895 15255 23905 15295
rect 23945 15255 23955 15295
rect 23995 15255 24005 15295
rect 24045 15255 24050 15295
rect 22850 15250 24050 15255
rect -1200 15195 0 15200
rect -1200 15155 -1195 15195
rect -1155 15155 -1145 15195
rect -1105 15155 -1095 15195
rect -1055 15155 -1045 15195
rect -1005 15155 -995 15195
rect -955 15155 0 15195
rect -1200 15150 0 15155
rect 22850 15195 24050 15200
rect 22850 15155 23805 15195
rect 23845 15155 23855 15195
rect 23895 15155 23905 15195
rect 23945 15155 23955 15195
rect 23995 15155 24005 15195
rect 24045 15155 24050 15195
rect 22850 15150 24050 15155
rect -1200 15095 0 15100
rect -1200 15055 -1195 15095
rect -1155 15055 -1145 15095
rect -1105 15055 -1095 15095
rect -1055 15055 -1045 15095
rect -1005 15055 -995 15095
rect -955 15055 0 15095
rect -1200 15050 0 15055
rect 22850 15095 24050 15100
rect 22850 15055 23805 15095
rect 23845 15055 23855 15095
rect 23895 15055 23905 15095
rect 23945 15055 23955 15095
rect 23995 15055 24005 15095
rect 24045 15055 24050 15095
rect 22850 15050 24050 15055
rect -1200 14995 0 15000
rect -1200 14955 -1195 14995
rect -1155 14955 -1145 14995
rect -1105 14955 -1095 14995
rect -1055 14955 -1045 14995
rect -1005 14955 -995 14995
rect -955 14955 0 14995
rect -1200 14950 0 14955
rect 22850 14995 24050 15000
rect 22850 14955 23805 14995
rect 23845 14955 23855 14995
rect 23895 14955 23905 14995
rect 23945 14955 23955 14995
rect 23995 14955 24005 14995
rect 24045 14955 24050 14995
rect 22850 14950 24050 14955
rect -1200 14895 0 14900
rect -1200 14855 -1195 14895
rect -1155 14855 -1145 14895
rect -1105 14855 -1095 14895
rect -1055 14855 -1045 14895
rect -1005 14855 -995 14895
rect -955 14855 0 14895
rect -1200 14850 0 14855
rect 22850 14895 24050 14900
rect 22850 14855 23805 14895
rect 23845 14855 23855 14895
rect 23895 14855 23905 14895
rect 23945 14855 23955 14895
rect 23995 14855 24005 14895
rect 24045 14855 24050 14895
rect 22850 14850 24050 14855
rect -1200 14795 0 14800
rect -1200 14755 -1195 14795
rect -1155 14755 -1145 14795
rect -1105 14755 -1095 14795
rect -1055 14755 -1045 14795
rect -1005 14755 -995 14795
rect -955 14755 0 14795
rect -1200 14750 0 14755
rect 22850 14795 24050 14800
rect 22850 14755 23805 14795
rect 23845 14755 23855 14795
rect 23895 14755 23905 14795
rect 23945 14755 23955 14795
rect 23995 14755 24005 14795
rect 24045 14755 24050 14795
rect 22850 14750 24050 14755
rect -1200 14695 0 14700
rect -1200 14655 -1195 14695
rect -1155 14655 -1145 14695
rect -1105 14655 -1095 14695
rect -1055 14655 -1045 14695
rect -1005 14655 -995 14695
rect -955 14655 0 14695
rect -1200 14650 0 14655
rect 22850 14695 24050 14700
rect 22850 14655 23805 14695
rect 23845 14655 23855 14695
rect 23895 14655 23905 14695
rect 23945 14655 23955 14695
rect 23995 14655 24005 14695
rect 24045 14655 24050 14695
rect 22850 14650 24050 14655
rect -900 14395 0 14400
rect -900 14355 -895 14395
rect -855 14355 -695 14395
rect -655 14355 -495 14395
rect -455 14355 -295 14395
rect -255 14355 -95 14395
rect -55 14355 0 14395
rect -900 14350 0 14355
rect 22850 14395 23750 14400
rect 22850 14355 22905 14395
rect 22945 14355 23305 14395
rect 23345 14355 23705 14395
rect 23745 14355 23750 14395
rect 22850 14350 23750 14355
rect 22250 14295 23650 14300
rect 22250 14255 23405 14295
rect 23445 14255 23455 14295
rect 23495 14255 23505 14295
rect 23545 14255 23555 14295
rect 23595 14255 23605 14295
rect 23645 14255 23650 14295
rect 22250 14245 23650 14255
rect 22250 14205 23405 14245
rect 23445 14205 23455 14245
rect 23495 14205 23505 14245
rect 23545 14205 23555 14245
rect 23595 14205 23605 14245
rect 23645 14205 23650 14245
rect 22250 14195 23650 14205
rect 22250 14155 23405 14195
rect 23445 14155 23455 14195
rect 23495 14155 23505 14195
rect 23545 14155 23555 14195
rect 23595 14155 23605 14195
rect 23645 14155 23650 14195
rect 22250 14145 23650 14155
rect 22250 14105 23405 14145
rect 23445 14105 23455 14145
rect 23495 14105 23505 14145
rect 23545 14105 23555 14145
rect 23595 14105 23605 14145
rect 23645 14105 23650 14145
rect 22250 14095 23650 14105
rect 22250 14055 23405 14095
rect 23445 14055 23455 14095
rect 23495 14055 23505 14095
rect 23545 14055 23555 14095
rect 23595 14055 23605 14095
rect 23645 14055 23650 14095
rect 22250 14050 23650 14055
rect -900 13995 0 14000
rect -900 13955 -895 13995
rect -855 13955 -695 13995
rect -655 13955 -495 13995
rect -455 13955 -295 13995
rect -255 13955 -95 13995
rect -55 13955 0 13995
rect -900 13950 0 13955
rect 22850 13995 23750 14000
rect 22850 13955 22905 13995
rect 22945 13955 23305 13995
rect 23345 13955 23705 13995
rect 23745 13955 23750 13995
rect 22850 13950 23750 13955
rect -900 13795 0 13800
rect -900 13755 -895 13795
rect -855 13755 -695 13795
rect -655 13755 -495 13795
rect -455 13755 -295 13795
rect -255 13755 -95 13795
rect -55 13755 0 13795
rect -900 13750 0 13755
rect -800 13695 600 13700
rect -800 13655 -795 13695
rect -755 13655 600 13695
rect -800 13650 600 13655
rect -900 13595 0 13600
rect -900 13555 -895 13595
rect -855 13555 -695 13595
rect -655 13555 -495 13595
rect -455 13555 -295 13595
rect -255 13555 -95 13595
rect -55 13555 0 13595
rect -900 13550 0 13555
rect 150 13495 200 13500
rect 150 13455 155 13495
rect 195 13455 200 13495
rect 150 13450 200 13455
rect 300 13495 350 13500
rect 300 13455 305 13495
rect 345 13455 350 13495
rect 300 13450 350 13455
rect -900 13395 0 13400
rect -900 13355 -895 13395
rect -855 13355 -695 13395
rect -655 13355 -495 13395
rect -455 13355 -295 13395
rect -255 13355 -95 13395
rect -55 13355 0 13395
rect -900 13350 0 13355
rect -600 13295 600 13300
rect -600 13255 -595 13295
rect -555 13255 600 13295
rect -600 13250 600 13255
rect -900 13195 0 13200
rect -900 13155 -895 13195
rect -855 13155 -695 13195
rect -655 13155 -495 13195
rect -455 13155 -295 13195
rect -255 13155 -95 13195
rect -55 13155 0 13195
rect -900 13150 0 13155
rect -900 12995 0 13000
rect -900 12955 -895 12995
rect -855 12955 -695 12995
rect -655 12955 -495 12995
rect -455 12955 -295 12995
rect -255 12955 -95 12995
rect -55 12955 0 12995
rect -900 12950 0 12955
rect 22850 12995 23750 13000
rect 22850 12955 22905 12995
rect 22945 12955 23305 12995
rect 23345 12955 23705 12995
rect 23745 12955 23750 12995
rect 22850 12950 23750 12955
rect 22250 12895 23250 12900
rect 22250 12855 23005 12895
rect 23045 12855 23055 12895
rect 23095 12855 23105 12895
rect 23145 12855 23155 12895
rect 23195 12855 23205 12895
rect 23245 12855 23250 12895
rect 22250 12845 23250 12855
rect 22250 12805 23005 12845
rect 23045 12805 23055 12845
rect 23095 12805 23105 12845
rect 23145 12805 23155 12845
rect 23195 12805 23205 12845
rect 23245 12805 23250 12845
rect 22250 12795 23250 12805
rect 22250 12755 23005 12795
rect 23045 12755 23055 12795
rect 23095 12755 23105 12795
rect 23145 12755 23155 12795
rect 23195 12755 23205 12795
rect 23245 12755 23250 12795
rect 22250 12745 23250 12755
rect 22250 12705 23005 12745
rect 23045 12705 23055 12745
rect 23095 12705 23105 12745
rect 23145 12705 23155 12745
rect 23195 12705 23205 12745
rect 23245 12705 23250 12745
rect 22250 12695 23250 12705
rect 22250 12655 23005 12695
rect 23045 12655 23055 12695
rect 23095 12655 23105 12695
rect 23145 12655 23155 12695
rect 23195 12655 23205 12695
rect 23245 12655 23250 12695
rect 22250 12650 23250 12655
rect -900 12595 0 12600
rect -900 12555 -895 12595
rect -855 12555 -695 12595
rect -655 12555 -495 12595
rect -455 12555 -295 12595
rect -255 12555 -95 12595
rect -55 12555 0 12595
rect -900 12550 0 12555
rect 22850 12595 23750 12600
rect 22850 12555 22905 12595
rect 22945 12555 23305 12595
rect 23345 12555 23705 12595
rect 23745 12555 23750 12595
rect 22850 12550 23750 12555
rect -1200 12295 0 12300
rect -1200 12255 -1195 12295
rect -1155 12255 -1145 12295
rect -1105 12255 -1095 12295
rect -1055 12255 -1045 12295
rect -1005 12255 -995 12295
rect -955 12255 0 12295
rect -1200 12250 0 12255
rect 22850 12295 24050 12300
rect 22850 12255 23805 12295
rect 23845 12255 23855 12295
rect 23895 12255 23905 12295
rect 23945 12255 23955 12295
rect 23995 12255 24005 12295
rect 24045 12255 24050 12295
rect 22850 12250 24050 12255
rect -1200 12195 0 12200
rect -1200 12155 -1195 12195
rect -1155 12155 -1145 12195
rect -1105 12155 -1095 12195
rect -1055 12155 -1045 12195
rect -1005 12155 -995 12195
rect -955 12155 0 12195
rect -1200 12150 0 12155
rect 22850 12195 24050 12200
rect 22850 12155 23805 12195
rect 23845 12155 23855 12195
rect 23895 12155 23905 12195
rect 23945 12155 23955 12195
rect 23995 12155 24005 12195
rect 24045 12155 24050 12195
rect 22850 12150 24050 12155
rect -1200 12095 0 12100
rect -1200 12055 -1195 12095
rect -1155 12055 -1145 12095
rect -1105 12055 -1095 12095
rect -1055 12055 -1045 12095
rect -1005 12055 -995 12095
rect -955 12055 0 12095
rect -1200 12050 0 12055
rect 22850 12095 24050 12100
rect 22850 12055 23805 12095
rect 23845 12055 23855 12095
rect 23895 12055 23905 12095
rect 23945 12055 23955 12095
rect 23995 12055 24005 12095
rect 24045 12055 24050 12095
rect 22850 12050 24050 12055
rect -1200 11995 0 12000
rect -1200 11955 -1195 11995
rect -1155 11955 -1145 11995
rect -1105 11955 -1095 11995
rect -1055 11955 -1045 11995
rect -1005 11955 -995 11995
rect -955 11955 0 11995
rect -1200 11950 0 11955
rect 22850 11995 24050 12000
rect 22850 11955 23805 11995
rect 23845 11955 23855 11995
rect 23895 11955 23905 11995
rect 23945 11955 23955 11995
rect 23995 11955 24005 11995
rect 24045 11955 24050 11995
rect 22850 11950 24050 11955
rect -1200 11895 0 11900
rect -1200 11855 -1195 11895
rect -1155 11855 -1145 11895
rect -1105 11855 -1095 11895
rect -1055 11855 -1045 11895
rect -1005 11855 -995 11895
rect -955 11855 0 11895
rect -1200 11850 0 11855
rect 22850 11895 24050 11900
rect 22850 11855 23805 11895
rect 23845 11855 23855 11895
rect 23895 11855 23905 11895
rect 23945 11855 23955 11895
rect 23995 11855 24005 11895
rect 24045 11855 24050 11895
rect 22850 11850 24050 11855
rect -1200 11795 0 11800
rect -1200 11755 -1195 11795
rect -1155 11755 -1145 11795
rect -1105 11755 -1095 11795
rect -1055 11755 -1045 11795
rect -1005 11755 -995 11795
rect -955 11755 0 11795
rect -1200 11750 0 11755
rect 22850 11795 24050 11800
rect 22850 11755 23805 11795
rect 23845 11755 23855 11795
rect 23895 11755 23905 11795
rect 23945 11755 23955 11795
rect 23995 11755 24005 11795
rect 24045 11755 24050 11795
rect 22850 11750 24050 11755
rect -1200 11695 0 11700
rect -1200 11655 -1195 11695
rect -1155 11655 -1145 11695
rect -1105 11655 -1095 11695
rect -1055 11655 -1045 11695
rect -1005 11655 -995 11695
rect -955 11655 0 11695
rect -1200 11650 0 11655
rect 22850 11695 24050 11700
rect 22850 11655 23805 11695
rect 23845 11655 23855 11695
rect 23895 11655 23905 11695
rect 23945 11655 23955 11695
rect 23995 11655 24005 11695
rect 24045 11655 24050 11695
rect 22850 11650 24050 11655
rect -1300 11595 24150 11600
rect -1300 11555 -1295 11595
rect -1255 11590 24105 11595
rect -1255 11560 10 11590
rect 40 11560 24105 11590
rect -1255 11555 24105 11560
rect 24145 11555 24150 11595
rect -1300 11545 24150 11555
rect -1300 11505 -1295 11545
rect -1255 11540 24105 11545
rect -1255 11510 10 11540
rect 40 11510 24105 11540
rect -1255 11505 24105 11510
rect 24145 11505 24150 11545
rect -1300 11500 24150 11505
rect -1200 11445 0 11450
rect -1200 11405 -1195 11445
rect -1155 11405 -1145 11445
rect -1105 11405 -1095 11445
rect -1055 11405 -1045 11445
rect -1005 11405 -995 11445
rect -955 11405 0 11445
rect -1200 11400 0 11405
rect 22850 11445 24050 11450
rect 22850 11405 23805 11445
rect 23845 11405 23855 11445
rect 23895 11405 23905 11445
rect 23945 11405 23955 11445
rect 23995 11405 24005 11445
rect 24045 11405 24050 11445
rect 22850 11400 24050 11405
rect -1200 11345 0 11350
rect -1200 11305 -1195 11345
rect -1155 11305 -1145 11345
rect -1105 11305 -1095 11345
rect -1055 11305 -1045 11345
rect -1005 11305 -995 11345
rect -955 11305 0 11345
rect -1200 11300 0 11305
rect 22850 11345 24050 11350
rect 22850 11305 23805 11345
rect 23845 11305 23855 11345
rect 23895 11305 23905 11345
rect 23945 11305 23955 11345
rect 23995 11305 24005 11345
rect 24045 11305 24050 11345
rect 22850 11300 24050 11305
rect -1200 11245 0 11250
rect -1200 11205 -1195 11245
rect -1155 11205 -1145 11245
rect -1105 11205 -1095 11245
rect -1055 11205 -1045 11245
rect -1005 11205 -995 11245
rect -955 11205 0 11245
rect -1200 11200 0 11205
rect 22850 11245 24050 11250
rect 22850 11205 23805 11245
rect 23845 11205 23855 11245
rect 23895 11205 23905 11245
rect 23945 11205 23955 11245
rect 23995 11205 24005 11245
rect 24045 11205 24050 11245
rect 22850 11200 24050 11205
rect -1200 11145 0 11150
rect -1200 11105 -1195 11145
rect -1155 11105 -1145 11145
rect -1105 11105 -1095 11145
rect -1055 11105 -1045 11145
rect -1005 11105 -995 11145
rect -955 11105 0 11145
rect -1200 11100 0 11105
rect 22850 11145 24050 11150
rect 22850 11105 23805 11145
rect 23845 11105 23855 11145
rect 23895 11105 23905 11145
rect 23945 11105 23955 11145
rect 23995 11105 24005 11145
rect 24045 11105 24050 11145
rect 22850 11100 24050 11105
rect -1200 11045 0 11050
rect -1200 11005 -1195 11045
rect -1155 11005 -1145 11045
rect -1105 11005 -1095 11045
rect -1055 11005 -1045 11045
rect -1005 11005 -995 11045
rect -955 11005 0 11045
rect -1200 11000 0 11005
rect 22850 11045 24050 11050
rect 22850 11005 23805 11045
rect 23845 11005 23855 11045
rect 23895 11005 23905 11045
rect 23945 11005 23955 11045
rect 23995 11005 24005 11045
rect 24045 11005 24050 11045
rect 22850 11000 24050 11005
rect -1200 10945 0 10950
rect -1200 10905 -1195 10945
rect -1155 10905 -1145 10945
rect -1105 10905 -1095 10945
rect -1055 10905 -1045 10945
rect -1005 10905 -995 10945
rect -955 10905 0 10945
rect -1200 10900 0 10905
rect 22850 10945 24050 10950
rect 22850 10905 23805 10945
rect 23845 10905 23855 10945
rect 23895 10905 23905 10945
rect 23945 10905 23955 10945
rect 23995 10905 24005 10945
rect 24045 10905 24050 10945
rect 22850 10900 24050 10905
rect -1200 10845 0 10850
rect -1200 10805 -1195 10845
rect -1155 10805 -1145 10845
rect -1105 10805 -1095 10845
rect -1055 10805 -1045 10845
rect -1005 10805 -995 10845
rect -955 10805 0 10845
rect -1200 10800 0 10805
rect 22850 10845 24050 10850
rect 22850 10805 23805 10845
rect 23845 10805 23855 10845
rect 23895 10805 23905 10845
rect 23945 10805 23955 10845
rect 23995 10805 24005 10845
rect 24045 10805 24050 10845
rect 22850 10800 24050 10805
rect -900 10545 0 10550
rect -900 10505 -895 10545
rect -855 10505 -695 10545
rect -655 10505 -495 10545
rect -455 10505 -295 10545
rect -255 10505 -95 10545
rect -55 10505 0 10545
rect -900 10500 0 10505
rect 22850 10545 23750 10550
rect 22850 10505 22905 10545
rect 22945 10505 23305 10545
rect 23345 10505 23705 10545
rect 23745 10505 23750 10545
rect 22850 10500 23750 10505
rect 22250 10445 23250 10450
rect 22250 10405 23005 10445
rect 23045 10405 23055 10445
rect 23095 10405 23105 10445
rect 23145 10405 23155 10445
rect 23195 10405 23205 10445
rect 23245 10405 23250 10445
rect 22250 10395 23250 10405
rect 22250 10355 23005 10395
rect 23045 10355 23055 10395
rect 23095 10355 23105 10395
rect 23145 10355 23155 10395
rect 23195 10355 23205 10395
rect 23245 10355 23250 10395
rect 22250 10345 23250 10355
rect 22250 10305 23005 10345
rect 23045 10305 23055 10345
rect 23095 10305 23105 10345
rect 23145 10305 23155 10345
rect 23195 10305 23205 10345
rect 23245 10305 23250 10345
rect 22250 10295 23250 10305
rect 22250 10255 23005 10295
rect 23045 10255 23055 10295
rect 23095 10255 23105 10295
rect 23145 10255 23155 10295
rect 23195 10255 23205 10295
rect 23245 10255 23250 10295
rect 22250 10245 23250 10255
rect 22250 10205 23005 10245
rect 23045 10205 23055 10245
rect 23095 10205 23105 10245
rect 23145 10205 23155 10245
rect 23195 10205 23205 10245
rect 23245 10205 23250 10245
rect 22250 10200 23250 10205
rect -900 10145 0 10150
rect -900 10105 -895 10145
rect -855 10105 -695 10145
rect -655 10105 -495 10145
rect -455 10105 -295 10145
rect -255 10105 -95 10145
rect -55 10105 0 10145
rect -900 10100 0 10105
rect 22850 10145 23750 10150
rect 22850 10105 22905 10145
rect 22945 10105 23305 10145
rect 23345 10105 23705 10145
rect 23745 10105 23750 10145
rect 22850 10100 23750 10105
rect -900 9945 0 9950
rect -900 9905 -895 9945
rect -855 9905 -695 9945
rect -655 9905 -495 9945
rect -455 9905 -295 9945
rect -255 9905 -95 9945
rect -55 9905 0 9945
rect -900 9900 0 9905
rect -200 9845 600 9850
rect -200 9805 -195 9845
rect -155 9805 600 9845
rect -200 9800 600 9805
rect -900 9745 0 9750
rect -900 9705 -895 9745
rect -855 9705 -695 9745
rect -655 9705 -495 9745
rect -455 9705 -295 9745
rect -255 9705 -95 9745
rect -55 9705 0 9745
rect -900 9700 0 9705
rect 150 9645 200 9650
rect 150 9605 155 9645
rect 195 9605 200 9645
rect 150 9600 200 9605
rect 300 9645 350 9650
rect 300 9605 305 9645
rect 345 9605 350 9645
rect 300 9600 350 9605
rect -900 9545 0 9550
rect -900 9505 -895 9545
rect -855 9505 -695 9545
rect -655 9505 -495 9545
rect -455 9505 -295 9545
rect -255 9505 -95 9545
rect -55 9505 0 9545
rect -900 9500 0 9505
rect -550 9400 -500 9450
rect -400 9445 600 9450
rect -400 9405 -395 9445
rect -355 9405 600 9445
rect -400 9400 600 9405
rect -900 9345 0 9350
rect -900 9305 -895 9345
rect -855 9305 -695 9345
rect -655 9305 -495 9345
rect -455 9305 -295 9345
rect -255 9305 -95 9345
rect -55 9305 0 9345
rect -900 9300 0 9305
rect -900 9145 0 9150
rect -900 9105 -895 9145
rect -855 9105 -695 9145
rect -655 9105 -495 9145
rect -455 9105 -295 9145
rect -255 9105 -95 9145
rect -55 9105 0 9145
rect -900 9100 0 9105
rect 22850 9145 23750 9150
rect 22850 9105 22905 9145
rect 22945 9105 23305 9145
rect 23345 9105 23705 9145
rect 23745 9105 23750 9145
rect 22850 9100 23750 9105
rect 22250 9045 23650 9050
rect 22250 9005 23405 9045
rect 23445 9005 23455 9045
rect 23495 9005 23505 9045
rect 23545 9005 23555 9045
rect 23595 9005 23605 9045
rect 23645 9005 23650 9045
rect 22250 8995 23650 9005
rect 22250 8955 23405 8995
rect 23445 8955 23455 8995
rect 23495 8955 23505 8995
rect 23545 8955 23555 8995
rect 23595 8955 23605 8995
rect 23645 8955 23650 8995
rect 22250 8945 23650 8955
rect 22250 8905 23405 8945
rect 23445 8905 23455 8945
rect 23495 8905 23505 8945
rect 23545 8905 23555 8945
rect 23595 8905 23605 8945
rect 23645 8905 23650 8945
rect 22250 8895 23650 8905
rect 22250 8855 23405 8895
rect 23445 8855 23455 8895
rect 23495 8855 23505 8895
rect 23545 8855 23555 8895
rect 23595 8855 23605 8895
rect 23645 8855 23650 8895
rect 22250 8845 23650 8855
rect 22250 8805 23405 8845
rect 23445 8805 23455 8845
rect 23495 8805 23505 8845
rect 23545 8805 23555 8845
rect 23595 8805 23605 8845
rect 23645 8805 23650 8845
rect 22250 8800 23650 8805
rect -900 8745 0 8750
rect -900 8705 -895 8745
rect -855 8705 -695 8745
rect -655 8705 -495 8745
rect -455 8705 -295 8745
rect -255 8705 -95 8745
rect -55 8705 0 8745
rect -900 8700 0 8705
rect 22850 8745 23750 8750
rect 22850 8705 22905 8745
rect 22945 8705 23305 8745
rect 23345 8705 23705 8745
rect 23745 8705 23750 8745
rect 22850 8700 23750 8705
rect -1200 8445 0 8450
rect -1200 8405 -1195 8445
rect -1155 8405 -1145 8445
rect -1105 8405 -1095 8445
rect -1055 8405 -1045 8445
rect -1005 8405 -995 8445
rect -955 8405 0 8445
rect -1200 8400 0 8405
rect 22850 8445 24050 8450
rect 22850 8405 23805 8445
rect 23845 8405 23855 8445
rect 23895 8405 23905 8445
rect 23945 8405 23955 8445
rect 23995 8405 24005 8445
rect 24045 8405 24050 8445
rect 22850 8400 24050 8405
rect -1200 8345 0 8350
rect -1200 8305 -1195 8345
rect -1155 8305 -1145 8345
rect -1105 8305 -1095 8345
rect -1055 8305 -1045 8345
rect -1005 8305 -995 8345
rect -955 8305 0 8345
rect -1200 8300 0 8305
rect 22850 8345 24050 8350
rect 22850 8305 23805 8345
rect 23845 8305 23855 8345
rect 23895 8305 23905 8345
rect 23945 8305 23955 8345
rect 23995 8305 24005 8345
rect 24045 8305 24050 8345
rect 22850 8300 24050 8305
rect -1200 8245 0 8250
rect -1200 8205 -1195 8245
rect -1155 8205 -1145 8245
rect -1105 8205 -1095 8245
rect -1055 8205 -1045 8245
rect -1005 8205 -995 8245
rect -955 8205 0 8245
rect -1200 8200 0 8205
rect 22850 8245 24050 8250
rect 22850 8205 23805 8245
rect 23845 8205 23855 8245
rect 23895 8205 23905 8245
rect 23945 8205 23955 8245
rect 23995 8205 24005 8245
rect 24045 8205 24050 8245
rect 22850 8200 24050 8205
rect -1200 8145 0 8150
rect -1200 8105 -1195 8145
rect -1155 8105 -1145 8145
rect -1105 8105 -1095 8145
rect -1055 8105 -1045 8145
rect -1005 8105 -995 8145
rect -955 8105 0 8145
rect -1200 8100 0 8105
rect 22850 8145 24050 8150
rect 22850 8105 23805 8145
rect 23845 8105 23855 8145
rect 23895 8105 23905 8145
rect 23945 8105 23955 8145
rect 23995 8105 24005 8145
rect 24045 8105 24050 8145
rect 22850 8100 24050 8105
rect -1200 8045 0 8050
rect -1200 8005 -1195 8045
rect -1155 8005 -1145 8045
rect -1105 8005 -1095 8045
rect -1055 8005 -1045 8045
rect -1005 8005 -995 8045
rect -955 8005 0 8045
rect -1200 8000 0 8005
rect 22850 8045 24050 8050
rect 22850 8005 23805 8045
rect 23845 8005 23855 8045
rect 23895 8005 23905 8045
rect 23945 8005 23955 8045
rect 23995 8005 24005 8045
rect 24045 8005 24050 8045
rect 22850 8000 24050 8005
rect -1200 7945 0 7950
rect -1200 7905 -1195 7945
rect -1155 7905 -1145 7945
rect -1105 7905 -1095 7945
rect -1055 7905 -1045 7945
rect -1005 7905 -995 7945
rect -955 7905 0 7945
rect -1200 7900 0 7905
rect 22850 7945 24050 7950
rect 22850 7905 23805 7945
rect 23845 7905 23855 7945
rect 23895 7905 23905 7945
rect 23945 7905 23955 7945
rect 23995 7905 24005 7945
rect 24045 7905 24050 7945
rect 22850 7900 24050 7905
rect -1200 7845 0 7850
rect -1200 7805 -1195 7845
rect -1155 7805 -1145 7845
rect -1105 7805 -1095 7845
rect -1055 7805 -1045 7845
rect -1005 7805 -995 7845
rect -955 7805 0 7845
rect -1200 7800 0 7805
rect 22850 7845 24050 7850
rect 22850 7805 23805 7845
rect 23845 7805 23855 7845
rect 23895 7805 23905 7845
rect 23945 7805 23955 7845
rect 23995 7805 24005 7845
rect 24045 7805 24050 7845
rect 22850 7800 24050 7805
<< via3 >>
rect -1195 15255 -1155 15295
rect -1145 15255 -1105 15295
rect -1095 15255 -1055 15295
rect -1045 15255 -1005 15295
rect -995 15255 -955 15295
rect 23805 15255 23845 15295
rect 23855 15255 23895 15295
rect 23905 15255 23945 15295
rect 23955 15255 23995 15295
rect 24005 15255 24045 15295
rect -1195 15155 -1155 15195
rect -1145 15155 -1105 15195
rect -1095 15155 -1055 15195
rect -1045 15155 -1005 15195
rect -995 15155 -955 15195
rect 23805 15155 23845 15195
rect 23855 15155 23895 15195
rect 23905 15155 23945 15195
rect 23955 15155 23995 15195
rect 24005 15155 24045 15195
rect -1195 15055 -1155 15095
rect -1145 15055 -1105 15095
rect -1095 15055 -1055 15095
rect -1045 15055 -1005 15095
rect -995 15055 -955 15095
rect 23805 15055 23845 15095
rect 23855 15055 23895 15095
rect 23905 15055 23945 15095
rect 23955 15055 23995 15095
rect 24005 15055 24045 15095
rect -1195 14955 -1155 14995
rect -1145 14955 -1105 14995
rect -1095 14955 -1055 14995
rect -1045 14955 -1005 14995
rect -995 14955 -955 14995
rect 23805 14955 23845 14995
rect 23855 14955 23895 14995
rect 23905 14955 23945 14995
rect 23955 14955 23995 14995
rect 24005 14955 24045 14995
rect -1195 14855 -1155 14895
rect -1145 14855 -1105 14895
rect -1095 14855 -1055 14895
rect -1045 14855 -1005 14895
rect -995 14855 -955 14895
rect 23805 14855 23845 14895
rect 23855 14855 23895 14895
rect 23905 14855 23945 14895
rect 23955 14855 23995 14895
rect 24005 14855 24045 14895
rect -1195 14755 -1155 14795
rect -1145 14755 -1105 14795
rect -1095 14755 -1055 14795
rect -1045 14755 -1005 14795
rect -995 14755 -955 14795
rect 23805 14755 23845 14795
rect 23855 14755 23895 14795
rect 23905 14755 23945 14795
rect 23955 14755 23995 14795
rect 24005 14755 24045 14795
rect -1195 14655 -1155 14695
rect -1145 14655 -1105 14695
rect -1095 14655 -1055 14695
rect -1045 14655 -1005 14695
rect -995 14655 -955 14695
rect 23805 14655 23845 14695
rect 23855 14655 23895 14695
rect 23905 14655 23945 14695
rect 23955 14655 23995 14695
rect 24005 14655 24045 14695
rect -895 14355 -855 14395
rect -695 14355 -655 14395
rect -495 14355 -455 14395
rect -295 14355 -255 14395
rect -95 14355 -55 14395
rect 22905 14355 22945 14395
rect 23305 14355 23345 14395
rect 23705 14355 23745 14395
rect 23405 14255 23445 14295
rect 23455 14255 23495 14295
rect 23505 14255 23545 14295
rect 23555 14255 23595 14295
rect 23605 14255 23645 14295
rect 23405 14205 23445 14245
rect 23455 14205 23495 14245
rect 23505 14205 23545 14245
rect 23555 14205 23595 14245
rect 23605 14205 23645 14245
rect 23405 14155 23445 14195
rect 23455 14155 23495 14195
rect 23505 14155 23545 14195
rect 23555 14155 23595 14195
rect 23605 14155 23645 14195
rect 23405 14105 23445 14145
rect 23455 14105 23495 14145
rect 23505 14105 23545 14145
rect 23555 14105 23595 14145
rect 23605 14105 23645 14145
rect 23405 14055 23445 14095
rect 23455 14055 23495 14095
rect 23505 14055 23545 14095
rect 23555 14055 23595 14095
rect 23605 14055 23645 14095
rect -895 13955 -855 13995
rect -695 13955 -655 13995
rect -495 13955 -455 13995
rect -295 13955 -255 13995
rect -95 13955 -55 13995
rect 22905 13955 22945 13995
rect 23305 13955 23345 13995
rect 23705 13955 23745 13995
rect -895 13755 -855 13795
rect -695 13755 -655 13795
rect -495 13755 -455 13795
rect -295 13755 -255 13795
rect -95 13755 -55 13795
rect -795 13655 -755 13695
rect -895 13555 -855 13595
rect -695 13555 -655 13595
rect -495 13555 -455 13595
rect -295 13555 -255 13595
rect -95 13555 -55 13595
rect 155 13490 195 13495
rect 155 13460 160 13490
rect 160 13460 190 13490
rect 190 13460 195 13490
rect 155 13455 195 13460
rect 305 13490 345 13495
rect 305 13460 310 13490
rect 310 13460 340 13490
rect 340 13460 345 13490
rect 305 13455 345 13460
rect -895 13355 -855 13395
rect -695 13355 -655 13395
rect -495 13355 -455 13395
rect -295 13355 -255 13395
rect -95 13355 -55 13395
rect -595 13255 -555 13295
rect -895 13155 -855 13195
rect -695 13155 -655 13195
rect -495 13155 -455 13195
rect -295 13155 -255 13195
rect -95 13155 -55 13195
rect -895 12955 -855 12995
rect -695 12955 -655 12995
rect -495 12955 -455 12995
rect -295 12955 -255 12995
rect -95 12955 -55 12995
rect 22905 12955 22945 12995
rect 23305 12955 23345 12995
rect 23705 12955 23745 12995
rect 23005 12855 23045 12895
rect 23055 12855 23095 12895
rect 23105 12855 23145 12895
rect 23155 12855 23195 12895
rect 23205 12855 23245 12895
rect 23005 12805 23045 12845
rect 23055 12805 23095 12845
rect 23105 12805 23145 12845
rect 23155 12805 23195 12845
rect 23205 12805 23245 12845
rect 23005 12755 23045 12795
rect 23055 12755 23095 12795
rect 23105 12755 23145 12795
rect 23155 12755 23195 12795
rect 23205 12755 23245 12795
rect 23005 12705 23045 12745
rect 23055 12705 23095 12745
rect 23105 12705 23145 12745
rect 23155 12705 23195 12745
rect 23205 12705 23245 12745
rect 23005 12655 23045 12695
rect 23055 12655 23095 12695
rect 23105 12655 23145 12695
rect 23155 12655 23195 12695
rect 23205 12655 23245 12695
rect -895 12555 -855 12595
rect -695 12555 -655 12595
rect -495 12555 -455 12595
rect -295 12555 -255 12595
rect -95 12555 -55 12595
rect 22905 12555 22945 12595
rect 23305 12555 23345 12595
rect 23705 12555 23745 12595
rect -1195 12255 -1155 12295
rect -1145 12255 -1105 12295
rect -1095 12255 -1055 12295
rect -1045 12255 -1005 12295
rect -995 12255 -955 12295
rect 23805 12255 23845 12295
rect 23855 12255 23895 12295
rect 23905 12255 23945 12295
rect 23955 12255 23995 12295
rect 24005 12255 24045 12295
rect -1195 12155 -1155 12195
rect -1145 12155 -1105 12195
rect -1095 12155 -1055 12195
rect -1045 12155 -1005 12195
rect -995 12155 -955 12195
rect 23805 12155 23845 12195
rect 23855 12155 23895 12195
rect 23905 12155 23945 12195
rect 23955 12155 23995 12195
rect 24005 12155 24045 12195
rect -1195 12055 -1155 12095
rect -1145 12055 -1105 12095
rect -1095 12055 -1055 12095
rect -1045 12055 -1005 12095
rect -995 12055 -955 12095
rect 23805 12055 23845 12095
rect 23855 12055 23895 12095
rect 23905 12055 23945 12095
rect 23955 12055 23995 12095
rect 24005 12055 24045 12095
rect -1195 11955 -1155 11995
rect -1145 11955 -1105 11995
rect -1095 11955 -1055 11995
rect -1045 11955 -1005 11995
rect -995 11955 -955 11995
rect 23805 11955 23845 11995
rect 23855 11955 23895 11995
rect 23905 11955 23945 11995
rect 23955 11955 23995 11995
rect 24005 11955 24045 11995
rect -1195 11855 -1155 11895
rect -1145 11855 -1105 11895
rect -1095 11855 -1055 11895
rect -1045 11855 -1005 11895
rect -995 11855 -955 11895
rect 23805 11855 23845 11895
rect 23855 11855 23895 11895
rect 23905 11855 23945 11895
rect 23955 11855 23995 11895
rect 24005 11855 24045 11895
rect -1195 11755 -1155 11795
rect -1145 11755 -1105 11795
rect -1095 11755 -1055 11795
rect -1045 11755 -1005 11795
rect -995 11755 -955 11795
rect 23805 11755 23845 11795
rect 23855 11755 23895 11795
rect 23905 11755 23945 11795
rect 23955 11755 23995 11795
rect 24005 11755 24045 11795
rect -1195 11655 -1155 11695
rect -1145 11655 -1105 11695
rect -1095 11655 -1055 11695
rect -1045 11655 -1005 11695
rect -995 11655 -955 11695
rect 23805 11655 23845 11695
rect 23855 11655 23895 11695
rect 23905 11655 23945 11695
rect 23955 11655 23995 11695
rect 24005 11655 24045 11695
rect -1295 11555 -1255 11595
rect 24105 11555 24145 11595
rect -1295 11505 -1255 11545
rect 24105 11505 24145 11545
rect -1195 11405 -1155 11445
rect -1145 11405 -1105 11445
rect -1095 11405 -1055 11445
rect -1045 11405 -1005 11445
rect -995 11405 -955 11445
rect 23805 11405 23845 11445
rect 23855 11405 23895 11445
rect 23905 11405 23945 11445
rect 23955 11405 23995 11445
rect 24005 11405 24045 11445
rect -1195 11305 -1155 11345
rect -1145 11305 -1105 11345
rect -1095 11305 -1055 11345
rect -1045 11305 -1005 11345
rect -995 11305 -955 11345
rect 23805 11305 23845 11345
rect 23855 11305 23895 11345
rect 23905 11305 23945 11345
rect 23955 11305 23995 11345
rect 24005 11305 24045 11345
rect -1195 11205 -1155 11245
rect -1145 11205 -1105 11245
rect -1095 11205 -1055 11245
rect -1045 11205 -1005 11245
rect -995 11205 -955 11245
rect 23805 11205 23845 11245
rect 23855 11205 23895 11245
rect 23905 11205 23945 11245
rect 23955 11205 23995 11245
rect 24005 11205 24045 11245
rect -1195 11105 -1155 11145
rect -1145 11105 -1105 11145
rect -1095 11105 -1055 11145
rect -1045 11105 -1005 11145
rect -995 11105 -955 11145
rect 23805 11105 23845 11145
rect 23855 11105 23895 11145
rect 23905 11105 23945 11145
rect 23955 11105 23995 11145
rect 24005 11105 24045 11145
rect -1195 11005 -1155 11045
rect -1145 11005 -1105 11045
rect -1095 11005 -1055 11045
rect -1045 11005 -1005 11045
rect -995 11005 -955 11045
rect 23805 11005 23845 11045
rect 23855 11005 23895 11045
rect 23905 11005 23945 11045
rect 23955 11005 23995 11045
rect 24005 11005 24045 11045
rect -1195 10905 -1155 10945
rect -1145 10905 -1105 10945
rect -1095 10905 -1055 10945
rect -1045 10905 -1005 10945
rect -995 10905 -955 10945
rect 23805 10905 23845 10945
rect 23855 10905 23895 10945
rect 23905 10905 23945 10945
rect 23955 10905 23995 10945
rect 24005 10905 24045 10945
rect -1195 10805 -1155 10845
rect -1145 10805 -1105 10845
rect -1095 10805 -1055 10845
rect -1045 10805 -1005 10845
rect -995 10805 -955 10845
rect 23805 10805 23845 10845
rect 23855 10805 23895 10845
rect 23905 10805 23945 10845
rect 23955 10805 23995 10845
rect 24005 10805 24045 10845
rect -895 10505 -855 10545
rect -695 10505 -655 10545
rect -495 10505 -455 10545
rect -295 10505 -255 10545
rect -95 10505 -55 10545
rect 22905 10505 22945 10545
rect 23305 10505 23345 10545
rect 23705 10505 23745 10545
rect 23005 10405 23045 10445
rect 23055 10405 23095 10445
rect 23105 10405 23145 10445
rect 23155 10405 23195 10445
rect 23205 10405 23245 10445
rect 23005 10355 23045 10395
rect 23055 10355 23095 10395
rect 23105 10355 23145 10395
rect 23155 10355 23195 10395
rect 23205 10355 23245 10395
rect 23005 10305 23045 10345
rect 23055 10305 23095 10345
rect 23105 10305 23145 10345
rect 23155 10305 23195 10345
rect 23205 10305 23245 10345
rect 23005 10255 23045 10295
rect 23055 10255 23095 10295
rect 23105 10255 23145 10295
rect 23155 10255 23195 10295
rect 23205 10255 23245 10295
rect 23005 10205 23045 10245
rect 23055 10205 23095 10245
rect 23105 10205 23145 10245
rect 23155 10205 23195 10245
rect 23205 10205 23245 10245
rect -895 10105 -855 10145
rect -695 10105 -655 10145
rect -495 10105 -455 10145
rect -295 10105 -255 10145
rect -95 10105 -55 10145
rect 22905 10105 22945 10145
rect 23305 10105 23345 10145
rect 23705 10105 23745 10145
rect -895 9905 -855 9945
rect -695 9905 -655 9945
rect -495 9905 -455 9945
rect -295 9905 -255 9945
rect -95 9905 -55 9945
rect -195 9805 -155 9845
rect -895 9705 -855 9745
rect -695 9705 -655 9745
rect -495 9705 -455 9745
rect -295 9705 -255 9745
rect -95 9705 -55 9745
rect 155 9640 195 9645
rect 155 9610 160 9640
rect 160 9610 190 9640
rect 190 9610 195 9640
rect 155 9605 195 9610
rect 305 9640 345 9645
rect 305 9610 310 9640
rect 310 9610 340 9640
rect 340 9610 345 9640
rect 305 9605 345 9610
rect -895 9505 -855 9545
rect -695 9505 -655 9545
rect -495 9505 -455 9545
rect -295 9505 -255 9545
rect -95 9505 -55 9545
rect -395 9405 -355 9445
rect -895 9305 -855 9345
rect -695 9305 -655 9345
rect -495 9305 -455 9345
rect -295 9305 -255 9345
rect -95 9305 -55 9345
rect -895 9105 -855 9145
rect -695 9105 -655 9145
rect -495 9105 -455 9145
rect -295 9105 -255 9145
rect -95 9105 -55 9145
rect 22905 9105 22945 9145
rect 23305 9105 23345 9145
rect 23705 9105 23745 9145
rect 23405 9005 23445 9045
rect 23455 9005 23495 9045
rect 23505 9005 23545 9045
rect 23555 9005 23595 9045
rect 23605 9005 23645 9045
rect 23405 8955 23445 8995
rect 23455 8955 23495 8995
rect 23505 8955 23545 8995
rect 23555 8955 23595 8995
rect 23605 8955 23645 8995
rect 23405 8905 23445 8945
rect 23455 8905 23495 8945
rect 23505 8905 23545 8945
rect 23555 8905 23595 8945
rect 23605 8905 23645 8945
rect 23405 8855 23445 8895
rect 23455 8855 23495 8895
rect 23505 8855 23545 8895
rect 23555 8855 23595 8895
rect 23605 8855 23645 8895
rect 23405 8805 23445 8845
rect 23455 8805 23495 8845
rect 23505 8805 23545 8845
rect 23555 8805 23595 8845
rect 23605 8805 23645 8845
rect -895 8705 -855 8745
rect -695 8705 -655 8745
rect -495 8705 -455 8745
rect -295 8705 -255 8745
rect -95 8705 -55 8745
rect 22905 8705 22945 8745
rect 23305 8705 23345 8745
rect 23705 8705 23745 8745
rect -1195 8405 -1155 8445
rect -1145 8405 -1105 8445
rect -1095 8405 -1055 8445
rect -1045 8405 -1005 8445
rect -995 8405 -955 8445
rect 23805 8405 23845 8445
rect 23855 8405 23895 8445
rect 23905 8405 23945 8445
rect 23955 8405 23995 8445
rect 24005 8405 24045 8445
rect -1195 8305 -1155 8345
rect -1145 8305 -1105 8345
rect -1095 8305 -1055 8345
rect -1045 8305 -1005 8345
rect -995 8305 -955 8345
rect 23805 8305 23845 8345
rect 23855 8305 23895 8345
rect 23905 8305 23945 8345
rect 23955 8305 23995 8345
rect 24005 8305 24045 8345
rect -1195 8205 -1155 8245
rect -1145 8205 -1105 8245
rect -1095 8205 -1055 8245
rect -1045 8205 -1005 8245
rect -995 8205 -955 8245
rect 23805 8205 23845 8245
rect 23855 8205 23895 8245
rect 23905 8205 23945 8245
rect 23955 8205 23995 8245
rect 24005 8205 24045 8245
rect -1195 8105 -1155 8145
rect -1145 8105 -1105 8145
rect -1095 8105 -1055 8145
rect -1045 8105 -1005 8145
rect -995 8105 -955 8145
rect 23805 8105 23845 8145
rect 23855 8105 23895 8145
rect 23905 8105 23945 8145
rect 23955 8105 23995 8145
rect 24005 8105 24045 8145
rect -1195 8005 -1155 8045
rect -1145 8005 -1105 8045
rect -1095 8005 -1055 8045
rect -1045 8005 -1005 8045
rect -995 8005 -955 8045
rect 23805 8005 23845 8045
rect 23855 8005 23895 8045
rect 23905 8005 23945 8045
rect 23955 8005 23995 8045
rect 24005 8005 24045 8045
rect -1195 7905 -1155 7945
rect -1145 7905 -1105 7945
rect -1095 7905 -1055 7945
rect -1045 7905 -1005 7945
rect -995 7905 -955 7945
rect 23805 7905 23845 7945
rect 23855 7905 23895 7945
rect 23905 7905 23945 7945
rect 23955 7905 23995 7945
rect 24005 7905 24045 7945
rect -1195 7805 -1155 7845
rect -1145 7805 -1105 7845
rect -1095 7805 -1055 7845
rect -1045 7805 -1005 7845
rect -995 7805 -955 7845
rect 23805 7805 23845 7845
rect 23855 7805 23895 7845
rect 23905 7805 23945 7845
rect 23955 7805 23995 7845
rect 24005 7805 24045 7845
<< metal4 >>
rect -1300 11595 -1250 15400
rect -1300 11555 -1295 11595
rect -1255 11555 -1250 11595
rect -1300 11545 -1250 11555
rect -1300 11505 -1295 11545
rect -1255 11505 -1250 11545
rect -1300 7700 -1250 11505
rect -1200 15295 -950 15400
rect -1200 15255 -1195 15295
rect -1155 15255 -1145 15295
rect -1105 15255 -1095 15295
rect -1055 15255 -1045 15295
rect -1005 15255 -995 15295
rect -955 15255 -950 15295
rect -1200 15195 -950 15255
rect -1200 15155 -1195 15195
rect -1155 15155 -1145 15195
rect -1105 15155 -1095 15195
rect -1055 15155 -1045 15195
rect -1005 15155 -995 15195
rect -955 15155 -950 15195
rect -1200 15095 -950 15155
rect -1200 15055 -1195 15095
rect -1155 15055 -1145 15095
rect -1105 15055 -1095 15095
rect -1055 15055 -1045 15095
rect -1005 15055 -995 15095
rect -955 15055 -950 15095
rect -1200 14995 -950 15055
rect -1200 14955 -1195 14995
rect -1155 14955 -1145 14995
rect -1105 14955 -1095 14995
rect -1055 14955 -1045 14995
rect -1005 14955 -995 14995
rect -955 14955 -950 14995
rect -1200 14895 -950 14955
rect -1200 14855 -1195 14895
rect -1155 14855 -1145 14895
rect -1105 14855 -1095 14895
rect -1055 14855 -1045 14895
rect -1005 14855 -995 14895
rect -955 14855 -950 14895
rect -1200 14795 -950 14855
rect -1200 14755 -1195 14795
rect -1155 14755 -1145 14795
rect -1105 14755 -1095 14795
rect -1055 14755 -1045 14795
rect -1005 14755 -995 14795
rect -955 14755 -950 14795
rect -1200 14695 -950 14755
rect -1200 14655 -1195 14695
rect -1155 14655 -1145 14695
rect -1105 14655 -1095 14695
rect -1055 14655 -1045 14695
rect -1005 14655 -995 14695
rect -955 14655 -950 14695
rect -1200 12295 -950 14655
rect -1200 12255 -1195 12295
rect -1155 12255 -1145 12295
rect -1105 12255 -1095 12295
rect -1055 12255 -1045 12295
rect -1005 12255 -995 12295
rect -955 12255 -950 12295
rect -1200 12195 -950 12255
rect -1200 12155 -1195 12195
rect -1155 12155 -1145 12195
rect -1105 12155 -1095 12195
rect -1055 12155 -1045 12195
rect -1005 12155 -995 12195
rect -955 12155 -950 12195
rect -1200 12095 -950 12155
rect -1200 12055 -1195 12095
rect -1155 12055 -1145 12095
rect -1105 12055 -1095 12095
rect -1055 12055 -1045 12095
rect -1005 12055 -995 12095
rect -955 12055 -950 12095
rect -1200 11995 -950 12055
rect -1200 11955 -1195 11995
rect -1155 11955 -1145 11995
rect -1105 11955 -1095 11995
rect -1055 11955 -1045 11995
rect -1005 11955 -995 11995
rect -955 11955 -950 11995
rect -1200 11895 -950 11955
rect -1200 11855 -1195 11895
rect -1155 11855 -1145 11895
rect -1105 11855 -1095 11895
rect -1055 11855 -1045 11895
rect -1005 11855 -995 11895
rect -955 11855 -950 11895
rect -1200 11795 -950 11855
rect -1200 11755 -1195 11795
rect -1155 11755 -1145 11795
rect -1105 11755 -1095 11795
rect -1055 11755 -1045 11795
rect -1005 11755 -995 11795
rect -955 11755 -950 11795
rect -1200 11695 -950 11755
rect -1200 11655 -1195 11695
rect -1155 11655 -1145 11695
rect -1105 11655 -1095 11695
rect -1055 11655 -1045 11695
rect -1005 11655 -995 11695
rect -955 11655 -950 11695
rect -1200 11445 -950 11655
rect -1200 11405 -1195 11445
rect -1155 11405 -1145 11445
rect -1105 11405 -1095 11445
rect -1055 11405 -1045 11445
rect -1005 11405 -995 11445
rect -955 11405 -950 11445
rect -1200 11345 -950 11405
rect -1200 11305 -1195 11345
rect -1155 11305 -1145 11345
rect -1105 11305 -1095 11345
rect -1055 11305 -1045 11345
rect -1005 11305 -995 11345
rect -955 11305 -950 11345
rect -1200 11245 -950 11305
rect -1200 11205 -1195 11245
rect -1155 11205 -1145 11245
rect -1105 11205 -1095 11245
rect -1055 11205 -1045 11245
rect -1005 11205 -995 11245
rect -955 11205 -950 11245
rect -1200 11145 -950 11205
rect -1200 11105 -1195 11145
rect -1155 11105 -1145 11145
rect -1105 11105 -1095 11145
rect -1055 11105 -1045 11145
rect -1005 11105 -995 11145
rect -955 11105 -950 11145
rect -1200 11045 -950 11105
rect -1200 11005 -1195 11045
rect -1155 11005 -1145 11045
rect -1105 11005 -1095 11045
rect -1055 11005 -1045 11045
rect -1005 11005 -995 11045
rect -955 11005 -950 11045
rect -1200 10945 -950 11005
rect -1200 10905 -1195 10945
rect -1155 10905 -1145 10945
rect -1105 10905 -1095 10945
rect -1055 10905 -1045 10945
rect -1005 10905 -995 10945
rect -955 10905 -950 10945
rect -1200 10845 -950 10905
rect -1200 10805 -1195 10845
rect -1155 10805 -1145 10845
rect -1105 10805 -1095 10845
rect -1055 10805 -1045 10845
rect -1005 10805 -995 10845
rect -955 10805 -950 10845
rect -1200 8445 -950 10805
rect -1200 8405 -1195 8445
rect -1155 8405 -1145 8445
rect -1105 8405 -1095 8445
rect -1055 8405 -1045 8445
rect -1005 8405 -995 8445
rect -955 8405 -950 8445
rect -1200 8345 -950 8405
rect -1200 8305 -1195 8345
rect -1155 8305 -1145 8345
rect -1105 8305 -1095 8345
rect -1055 8305 -1045 8345
rect -1005 8305 -995 8345
rect -955 8305 -950 8345
rect -1200 8245 -950 8305
rect -1200 8205 -1195 8245
rect -1155 8205 -1145 8245
rect -1105 8205 -1095 8245
rect -1055 8205 -1045 8245
rect -1005 8205 -995 8245
rect -955 8205 -950 8245
rect -1200 8145 -950 8205
rect -1200 8105 -1195 8145
rect -1155 8105 -1145 8145
rect -1105 8105 -1095 8145
rect -1055 8105 -1045 8145
rect -1005 8105 -995 8145
rect -955 8105 -950 8145
rect -1200 8045 -950 8105
rect -1200 8005 -1195 8045
rect -1155 8005 -1145 8045
rect -1105 8005 -1095 8045
rect -1055 8005 -1045 8045
rect -1005 8005 -995 8045
rect -955 8005 -950 8045
rect -1200 7945 -950 8005
rect -1200 7905 -1195 7945
rect -1155 7905 -1145 7945
rect -1105 7905 -1095 7945
rect -1055 7905 -1045 7945
rect -1005 7905 -995 7945
rect -955 7905 -950 7945
rect -1200 7845 -950 7905
rect -1200 7805 -1195 7845
rect -1155 7805 -1145 7845
rect -1105 7805 -1095 7845
rect -1055 7805 -1045 7845
rect -1005 7805 -995 7845
rect -955 7805 -950 7845
rect -1200 7700 -950 7805
rect -900 14395 -850 15400
rect -900 14355 -895 14395
rect -855 14355 -850 14395
rect -900 13995 -850 14355
rect -900 13955 -895 13995
rect -855 13955 -850 13995
rect -900 13795 -850 13955
rect -900 13755 -895 13795
rect -855 13755 -850 13795
rect -900 13595 -850 13755
rect -900 13555 -895 13595
rect -855 13555 -850 13595
rect -900 13395 -850 13555
rect -900 13355 -895 13395
rect -855 13355 -850 13395
rect -900 13195 -850 13355
rect -900 13155 -895 13195
rect -855 13155 -850 13195
rect -900 12995 -850 13155
rect -900 12955 -895 12995
rect -855 12955 -850 12995
rect -900 12595 -850 12955
rect -900 12555 -895 12595
rect -855 12555 -850 12595
rect -900 10545 -850 12555
rect -900 10505 -895 10545
rect -855 10505 -850 10545
rect -900 10145 -850 10505
rect -900 10105 -895 10145
rect -855 10105 -850 10145
rect -900 9945 -850 10105
rect -900 9905 -895 9945
rect -855 9905 -850 9945
rect -900 9745 -850 9905
rect -900 9705 -895 9745
rect -855 9705 -850 9745
rect -900 9545 -850 9705
rect -900 9505 -895 9545
rect -855 9505 -850 9545
rect -900 9345 -850 9505
rect -900 9305 -895 9345
rect -855 9305 -850 9345
rect -900 9145 -850 9305
rect -900 9105 -895 9145
rect -855 9105 -850 9145
rect -900 8745 -850 9105
rect -900 8705 -895 8745
rect -855 8705 -850 8745
rect -900 7700 -850 8705
rect -800 13695 -750 15400
rect -800 13655 -795 13695
rect -755 13655 -750 13695
rect -800 7700 -750 13655
rect -700 14395 -650 15400
rect -700 14355 -695 14395
rect -655 14355 -650 14395
rect -700 13995 -650 14355
rect -700 13955 -695 13995
rect -655 13955 -650 13995
rect -700 13795 -650 13955
rect -700 13755 -695 13795
rect -655 13755 -650 13795
rect -700 13595 -650 13755
rect -700 13555 -695 13595
rect -655 13555 -650 13595
rect -700 13395 -650 13555
rect -700 13355 -695 13395
rect -655 13355 -650 13395
rect -700 13195 -650 13355
rect -700 13155 -695 13195
rect -655 13155 -650 13195
rect -700 12995 -650 13155
rect -700 12955 -695 12995
rect -655 12955 -650 12995
rect -700 12595 -650 12955
rect -700 12555 -695 12595
rect -655 12555 -650 12595
rect -700 10545 -650 12555
rect -700 10505 -695 10545
rect -655 10505 -650 10545
rect -700 10145 -650 10505
rect -700 10105 -695 10145
rect -655 10105 -650 10145
rect -700 9945 -650 10105
rect -700 9905 -695 9945
rect -655 9905 -650 9945
rect -700 9745 -650 9905
rect -700 9705 -695 9745
rect -655 9705 -650 9745
rect -700 9545 -650 9705
rect -700 9505 -695 9545
rect -655 9505 -650 9545
rect -700 9345 -650 9505
rect -700 9305 -695 9345
rect -655 9305 -650 9345
rect -700 9145 -650 9305
rect -700 9105 -695 9145
rect -655 9105 -650 9145
rect -700 8745 -650 9105
rect -700 8705 -695 8745
rect -655 8705 -650 8745
rect -700 7700 -650 8705
rect -600 13295 -550 15400
rect -600 13255 -595 13295
rect -555 13255 -550 13295
rect -600 7700 -550 13255
rect -500 14395 -450 15400
rect -500 14355 -495 14395
rect -455 14355 -450 14395
rect -500 13995 -450 14355
rect -500 13955 -495 13995
rect -455 13955 -450 13995
rect -500 13795 -450 13955
rect -500 13755 -495 13795
rect -455 13755 -450 13795
rect -500 13595 -450 13755
rect -500 13555 -495 13595
rect -455 13555 -450 13595
rect -500 13395 -450 13555
rect -500 13355 -495 13395
rect -455 13355 -450 13395
rect -500 13195 -450 13355
rect -500 13155 -495 13195
rect -455 13155 -450 13195
rect -500 12995 -450 13155
rect -500 12955 -495 12995
rect -455 12955 -450 12995
rect -500 12595 -450 12955
rect -500 12555 -495 12595
rect -455 12555 -450 12595
rect -500 10545 -450 12555
rect -500 10505 -495 10545
rect -455 10505 -450 10545
rect -500 10145 -450 10505
rect -500 10105 -495 10145
rect -455 10105 -450 10145
rect -500 9945 -450 10105
rect -500 9905 -495 9945
rect -455 9905 -450 9945
rect -500 9745 -450 9905
rect -500 9705 -495 9745
rect -455 9705 -450 9745
rect -500 9545 -450 9705
rect -500 9505 -495 9545
rect -455 9505 -450 9545
rect -500 9345 -450 9505
rect -500 9305 -495 9345
rect -455 9305 -450 9345
rect -500 9145 -450 9305
rect -500 9105 -495 9145
rect -455 9105 -450 9145
rect -500 8745 -450 9105
rect -500 8705 -495 8745
rect -455 8705 -450 8745
rect -500 7700 -450 8705
rect -400 9445 -350 15400
rect -400 9405 -395 9445
rect -355 9405 -350 9445
rect -400 7700 -350 9405
rect -300 14395 -250 15400
rect -300 14355 -295 14395
rect -255 14355 -250 14395
rect -300 13995 -250 14355
rect -300 13955 -295 13995
rect -255 13955 -250 13995
rect -300 13795 -250 13955
rect -300 13755 -295 13795
rect -255 13755 -250 13795
rect -300 13595 -250 13755
rect -300 13555 -295 13595
rect -255 13555 -250 13595
rect -300 13395 -250 13555
rect -300 13355 -295 13395
rect -255 13355 -250 13395
rect -300 13195 -250 13355
rect -300 13155 -295 13195
rect -255 13155 -250 13195
rect -300 12995 -250 13155
rect -300 12955 -295 12995
rect -255 12955 -250 12995
rect -300 12595 -250 12955
rect -300 12555 -295 12595
rect -255 12555 -250 12595
rect -300 10545 -250 12555
rect -300 10505 -295 10545
rect -255 10505 -250 10545
rect -300 10145 -250 10505
rect -300 10105 -295 10145
rect -255 10105 -250 10145
rect -300 9945 -250 10105
rect -300 9905 -295 9945
rect -255 9905 -250 9945
rect -300 9745 -250 9905
rect -300 9705 -295 9745
rect -255 9705 -250 9745
rect -300 9545 -250 9705
rect -300 9505 -295 9545
rect -255 9505 -250 9545
rect -300 9345 -250 9505
rect -300 9305 -295 9345
rect -255 9305 -250 9345
rect -300 9145 -250 9305
rect -300 9105 -295 9145
rect -255 9105 -250 9145
rect -300 8745 -250 9105
rect -300 8705 -295 8745
rect -255 8705 -250 8745
rect -300 7700 -250 8705
rect -200 9845 -150 15400
rect -200 9805 -195 9845
rect -155 9805 -150 9845
rect -200 9250 -150 9805
rect -100 14395 -50 15400
rect -100 14355 -95 14395
rect -55 14355 -50 14395
rect -100 13995 -50 14355
rect -100 13955 -95 13995
rect -55 13955 -50 13995
rect -100 13795 -50 13955
rect -100 13755 -95 13795
rect -55 13755 -50 13795
rect -100 13595 -50 13755
rect -100 13555 -95 13595
rect -55 13555 -50 13595
rect -100 13395 -50 13555
rect -100 13355 -95 13395
rect -55 13355 -50 13395
rect -100 13195 -50 13355
rect -100 13155 -95 13195
rect -55 13155 -50 13195
rect -100 12995 -50 13155
rect -100 12955 -95 12995
rect -55 12955 -50 12995
rect -100 12595 -50 12955
rect -100 12555 -95 12595
rect -55 12555 -50 12595
rect -100 10545 -50 12555
rect -100 10505 -95 10545
rect -55 10505 -50 10545
rect -100 10145 -50 10505
rect -100 10105 -95 10145
rect -55 10105 -50 10145
rect -100 9945 -50 10105
rect -100 9905 -95 9945
rect -55 9905 -50 9945
rect -100 9745 -50 9905
rect -100 9705 -95 9745
rect -55 9705 -50 9745
rect -100 9545 -50 9705
rect -100 9505 -95 9545
rect -55 9505 -50 9545
rect -100 9345 -50 9505
rect -100 9305 -95 9345
rect -55 9305 -50 9345
rect -200 9200 -155 9250
rect -200 7700 -150 9200
rect -100 9145 -50 9305
rect 150 13495 200 15400
rect 150 13455 155 13495
rect 195 13455 200 13495
rect 150 9645 200 13455
rect 150 9605 155 9645
rect 195 9605 200 9645
rect 150 9250 200 9605
rect 149 9199 200 9250
rect -100 9105 -95 9145
rect -55 9105 -50 9145
rect -100 8745 -50 9105
rect -100 8705 -95 8745
rect -55 8705 -50 8745
rect -100 7700 -50 8705
rect 150 7700 200 9199
rect 300 13495 350 15400
rect 300 13455 305 13495
rect 345 13455 350 13495
rect 300 9645 350 13455
rect 300 9605 305 9645
rect 345 9605 350 9645
rect 300 9251 350 9605
rect 22900 14395 22950 15400
rect 22900 14355 22905 14395
rect 22945 14355 22950 14395
rect 22900 13995 22950 14355
rect 22900 13955 22905 13995
rect 22945 13955 22950 13995
rect 22900 12995 22950 13955
rect 22900 12955 22905 12995
rect 22945 12955 22950 12995
rect 22900 12595 22950 12955
rect 22900 12555 22905 12595
rect 22945 12555 22950 12595
rect 22900 10545 22950 12555
rect 22900 10505 22905 10545
rect 22945 10505 22950 10545
rect 22900 10145 22950 10505
rect 22900 10105 22905 10145
rect 22945 10105 22950 10145
rect 300 9200 351 9251
rect 300 7700 350 9200
rect 22900 9145 22950 10105
rect 22900 9105 22905 9145
rect 22945 9105 22950 9145
rect 22900 8745 22950 9105
rect 22900 8705 22905 8745
rect 22945 8705 22950 8745
rect 22900 7700 22950 8705
rect 23000 12895 23250 15400
rect 23000 12855 23005 12895
rect 23045 12855 23055 12895
rect 23095 12855 23105 12895
rect 23145 12855 23155 12895
rect 23195 12855 23205 12895
rect 23245 12855 23250 12895
rect 23000 12845 23250 12855
rect 23000 12805 23005 12845
rect 23045 12805 23055 12845
rect 23095 12805 23105 12845
rect 23145 12805 23155 12845
rect 23195 12805 23205 12845
rect 23245 12805 23250 12845
rect 23000 12795 23250 12805
rect 23000 12755 23005 12795
rect 23045 12755 23055 12795
rect 23095 12755 23105 12795
rect 23145 12755 23155 12795
rect 23195 12755 23205 12795
rect 23245 12755 23250 12795
rect 23000 12745 23250 12755
rect 23000 12705 23005 12745
rect 23045 12705 23055 12745
rect 23095 12705 23105 12745
rect 23145 12705 23155 12745
rect 23195 12705 23205 12745
rect 23245 12705 23250 12745
rect 23000 12695 23250 12705
rect 23000 12655 23005 12695
rect 23045 12655 23055 12695
rect 23095 12655 23105 12695
rect 23145 12655 23155 12695
rect 23195 12655 23205 12695
rect 23245 12655 23250 12695
rect 23000 10445 23250 12655
rect 23000 10405 23005 10445
rect 23045 10405 23055 10445
rect 23095 10405 23105 10445
rect 23145 10405 23155 10445
rect 23195 10405 23205 10445
rect 23245 10405 23250 10445
rect 23000 10395 23250 10405
rect 23000 10355 23005 10395
rect 23045 10355 23055 10395
rect 23095 10355 23105 10395
rect 23145 10355 23155 10395
rect 23195 10355 23205 10395
rect 23245 10355 23250 10395
rect 23000 10345 23250 10355
rect 23000 10305 23005 10345
rect 23045 10305 23055 10345
rect 23095 10305 23105 10345
rect 23145 10305 23155 10345
rect 23195 10305 23205 10345
rect 23245 10305 23250 10345
rect 23000 10295 23250 10305
rect 23000 10255 23005 10295
rect 23045 10255 23055 10295
rect 23095 10255 23105 10295
rect 23145 10255 23155 10295
rect 23195 10255 23205 10295
rect 23245 10255 23250 10295
rect 23000 10245 23250 10255
rect 23000 10205 23005 10245
rect 23045 10205 23055 10245
rect 23095 10205 23105 10245
rect 23145 10205 23155 10245
rect 23195 10205 23205 10245
rect 23245 10205 23250 10245
rect 23000 7700 23250 10205
rect 23300 14395 23350 15400
rect 23300 14355 23305 14395
rect 23345 14355 23350 14395
rect 23300 13995 23350 14355
rect 23300 13955 23305 13995
rect 23345 13955 23350 13995
rect 23300 12995 23350 13955
rect 23300 12955 23305 12995
rect 23345 12955 23350 12995
rect 23300 12595 23350 12955
rect 23300 12555 23305 12595
rect 23345 12555 23350 12595
rect 23300 10545 23350 12555
rect 23300 10505 23305 10545
rect 23345 10505 23350 10545
rect 23300 10145 23350 10505
rect 23300 10105 23305 10145
rect 23345 10105 23350 10145
rect 23300 9145 23350 10105
rect 23300 9105 23305 9145
rect 23345 9105 23350 9145
rect 23300 8745 23350 9105
rect 23300 8705 23305 8745
rect 23345 8705 23350 8745
rect 23300 7700 23350 8705
rect 23400 14295 23650 15400
rect 23400 14255 23405 14295
rect 23445 14255 23455 14295
rect 23495 14255 23505 14295
rect 23545 14255 23555 14295
rect 23595 14255 23605 14295
rect 23645 14255 23650 14295
rect 23400 14245 23650 14255
rect 23400 14205 23405 14245
rect 23445 14205 23455 14245
rect 23495 14205 23505 14245
rect 23545 14205 23555 14245
rect 23595 14205 23605 14245
rect 23645 14205 23650 14245
rect 23400 14195 23650 14205
rect 23400 14155 23405 14195
rect 23445 14155 23455 14195
rect 23495 14155 23505 14195
rect 23545 14155 23555 14195
rect 23595 14155 23605 14195
rect 23645 14155 23650 14195
rect 23400 14145 23650 14155
rect 23400 14105 23405 14145
rect 23445 14105 23455 14145
rect 23495 14105 23505 14145
rect 23545 14105 23555 14145
rect 23595 14105 23605 14145
rect 23645 14105 23650 14145
rect 23400 14095 23650 14105
rect 23400 14055 23405 14095
rect 23445 14055 23455 14095
rect 23495 14055 23505 14095
rect 23545 14055 23555 14095
rect 23595 14055 23605 14095
rect 23645 14055 23650 14095
rect 23400 9045 23650 14055
rect 23400 9005 23405 9045
rect 23445 9005 23455 9045
rect 23495 9005 23505 9045
rect 23545 9005 23555 9045
rect 23595 9005 23605 9045
rect 23645 9005 23650 9045
rect 23400 8995 23650 9005
rect 23400 8955 23405 8995
rect 23445 8955 23455 8995
rect 23495 8955 23505 8995
rect 23545 8955 23555 8995
rect 23595 8955 23605 8995
rect 23645 8955 23650 8995
rect 23400 8945 23650 8955
rect 23400 8905 23405 8945
rect 23445 8905 23455 8945
rect 23495 8905 23505 8945
rect 23545 8905 23555 8945
rect 23595 8905 23605 8945
rect 23645 8905 23650 8945
rect 23400 8895 23650 8905
rect 23400 8855 23405 8895
rect 23445 8855 23455 8895
rect 23495 8855 23505 8895
rect 23545 8855 23555 8895
rect 23595 8855 23605 8895
rect 23645 8855 23650 8895
rect 23400 8845 23650 8855
rect 23400 8805 23405 8845
rect 23445 8805 23455 8845
rect 23495 8805 23505 8845
rect 23545 8805 23555 8845
rect 23595 8805 23605 8845
rect 23645 8805 23650 8845
rect 23400 7700 23650 8805
rect 23700 14395 23750 15400
rect 23700 14355 23705 14395
rect 23745 14355 23750 14395
rect 23700 13995 23750 14355
rect 23700 13955 23705 13995
rect 23745 13955 23750 13995
rect 23700 12995 23750 13955
rect 23700 12955 23705 12995
rect 23745 12955 23750 12995
rect 23700 12595 23750 12955
rect 23700 12555 23705 12595
rect 23745 12555 23750 12595
rect 23700 10545 23750 12555
rect 23700 10505 23705 10545
rect 23745 10505 23750 10545
rect 23700 10145 23750 10505
rect 23700 10105 23705 10145
rect 23745 10105 23750 10145
rect 23700 9145 23750 10105
rect 23700 9105 23705 9145
rect 23745 9105 23750 9145
rect 23700 8745 23750 9105
rect 23700 8705 23705 8745
rect 23745 8705 23750 8745
rect 23700 7700 23750 8705
rect 23800 15295 24050 15400
rect 23800 15255 23805 15295
rect 23845 15255 23855 15295
rect 23895 15255 23905 15295
rect 23945 15255 23955 15295
rect 23995 15255 24005 15295
rect 24045 15255 24050 15295
rect 23800 15195 24050 15255
rect 23800 15155 23805 15195
rect 23845 15155 23855 15195
rect 23895 15155 23905 15195
rect 23945 15155 23955 15195
rect 23995 15155 24005 15195
rect 24045 15155 24050 15195
rect 23800 15095 24050 15155
rect 23800 15055 23805 15095
rect 23845 15055 23855 15095
rect 23895 15055 23905 15095
rect 23945 15055 23955 15095
rect 23995 15055 24005 15095
rect 24045 15055 24050 15095
rect 23800 14995 24050 15055
rect 23800 14955 23805 14995
rect 23845 14955 23855 14995
rect 23895 14955 23905 14995
rect 23945 14955 23955 14995
rect 23995 14955 24005 14995
rect 24045 14955 24050 14995
rect 23800 14895 24050 14955
rect 23800 14855 23805 14895
rect 23845 14855 23855 14895
rect 23895 14855 23905 14895
rect 23945 14855 23955 14895
rect 23995 14855 24005 14895
rect 24045 14855 24050 14895
rect 23800 14795 24050 14855
rect 23800 14755 23805 14795
rect 23845 14755 23855 14795
rect 23895 14755 23905 14795
rect 23945 14755 23955 14795
rect 23995 14755 24005 14795
rect 24045 14755 24050 14795
rect 23800 14695 24050 14755
rect 23800 14655 23805 14695
rect 23845 14655 23855 14695
rect 23895 14655 23905 14695
rect 23945 14655 23955 14695
rect 23995 14655 24005 14695
rect 24045 14655 24050 14695
rect 23800 12295 24050 14655
rect 23800 12255 23805 12295
rect 23845 12255 23855 12295
rect 23895 12255 23905 12295
rect 23945 12255 23955 12295
rect 23995 12255 24005 12295
rect 24045 12255 24050 12295
rect 23800 12195 24050 12255
rect 23800 12155 23805 12195
rect 23845 12155 23855 12195
rect 23895 12155 23905 12195
rect 23945 12155 23955 12195
rect 23995 12155 24005 12195
rect 24045 12155 24050 12195
rect 23800 12095 24050 12155
rect 23800 12055 23805 12095
rect 23845 12055 23855 12095
rect 23895 12055 23905 12095
rect 23945 12055 23955 12095
rect 23995 12055 24005 12095
rect 24045 12055 24050 12095
rect 23800 11995 24050 12055
rect 23800 11955 23805 11995
rect 23845 11955 23855 11995
rect 23895 11955 23905 11995
rect 23945 11955 23955 11995
rect 23995 11955 24005 11995
rect 24045 11955 24050 11995
rect 23800 11895 24050 11955
rect 23800 11855 23805 11895
rect 23845 11855 23855 11895
rect 23895 11855 23905 11895
rect 23945 11855 23955 11895
rect 23995 11855 24005 11895
rect 24045 11855 24050 11895
rect 23800 11795 24050 11855
rect 23800 11755 23805 11795
rect 23845 11755 23855 11795
rect 23895 11755 23905 11795
rect 23945 11755 23955 11795
rect 23995 11755 24005 11795
rect 24045 11755 24050 11795
rect 23800 11695 24050 11755
rect 23800 11655 23805 11695
rect 23845 11655 23855 11695
rect 23895 11655 23905 11695
rect 23945 11655 23955 11695
rect 23995 11655 24005 11695
rect 24045 11655 24050 11695
rect 23800 11445 24050 11655
rect 23800 11405 23805 11445
rect 23845 11405 23855 11445
rect 23895 11405 23905 11445
rect 23945 11405 23955 11445
rect 23995 11405 24005 11445
rect 24045 11405 24050 11445
rect 23800 11345 24050 11405
rect 23800 11305 23805 11345
rect 23845 11305 23855 11345
rect 23895 11305 23905 11345
rect 23945 11305 23955 11345
rect 23995 11305 24005 11345
rect 24045 11305 24050 11345
rect 23800 11245 24050 11305
rect 23800 11205 23805 11245
rect 23845 11205 23855 11245
rect 23895 11205 23905 11245
rect 23945 11205 23955 11245
rect 23995 11205 24005 11245
rect 24045 11205 24050 11245
rect 23800 11145 24050 11205
rect 23800 11105 23805 11145
rect 23845 11105 23855 11145
rect 23895 11105 23905 11145
rect 23945 11105 23955 11145
rect 23995 11105 24005 11145
rect 24045 11105 24050 11145
rect 23800 11045 24050 11105
rect 23800 11005 23805 11045
rect 23845 11005 23855 11045
rect 23895 11005 23905 11045
rect 23945 11005 23955 11045
rect 23995 11005 24005 11045
rect 24045 11005 24050 11045
rect 23800 10945 24050 11005
rect 23800 10905 23805 10945
rect 23845 10905 23855 10945
rect 23895 10905 23905 10945
rect 23945 10905 23955 10945
rect 23995 10905 24005 10945
rect 24045 10905 24050 10945
rect 23800 10845 24050 10905
rect 23800 10805 23805 10845
rect 23845 10805 23855 10845
rect 23895 10805 23905 10845
rect 23945 10805 23955 10845
rect 23995 10805 24005 10845
rect 24045 10805 24050 10845
rect 23800 8445 24050 10805
rect 23800 8405 23805 8445
rect 23845 8405 23855 8445
rect 23895 8405 23905 8445
rect 23945 8405 23955 8445
rect 23995 8405 24005 8445
rect 24045 8405 24050 8445
rect 23800 8345 24050 8405
rect 23800 8305 23805 8345
rect 23845 8305 23855 8345
rect 23895 8305 23905 8345
rect 23945 8305 23955 8345
rect 23995 8305 24005 8345
rect 24045 8305 24050 8345
rect 23800 8245 24050 8305
rect 23800 8205 23805 8245
rect 23845 8205 23855 8245
rect 23895 8205 23905 8245
rect 23945 8205 23955 8245
rect 23995 8205 24005 8245
rect 24045 8205 24050 8245
rect 23800 8145 24050 8205
rect 23800 8105 23805 8145
rect 23845 8105 23855 8145
rect 23895 8105 23905 8145
rect 23945 8105 23955 8145
rect 23995 8105 24005 8145
rect 24045 8105 24050 8145
rect 23800 8045 24050 8105
rect 23800 8005 23805 8045
rect 23845 8005 23855 8045
rect 23895 8005 23905 8045
rect 23945 8005 23955 8045
rect 23995 8005 24005 8045
rect 24045 8005 24050 8045
rect 23800 7945 24050 8005
rect 23800 7905 23805 7945
rect 23845 7905 23855 7945
rect 23895 7905 23905 7945
rect 23945 7905 23955 7945
rect 23995 7905 24005 7945
rect 24045 7905 24050 7945
rect 23800 7845 24050 7905
rect 23800 7805 23805 7845
rect 23845 7805 23855 7845
rect 23895 7805 23905 7845
rect 23945 7805 23955 7845
rect 23995 7805 24005 7845
rect 24045 7805 24050 7845
rect 23800 7700 24050 7805
rect 24100 11595 24150 15400
rect 24100 11555 24105 11595
rect 24145 11555 24150 11595
rect 24100 11545 24150 11555
rect 24100 11505 24105 11545
rect 24145 11505 24150 11545
rect 24100 7700 24150 11505
use ddaa_slice  ddaa_slice_0
timestamp 1726841226
transform 1 0 550 0 1 11550
box 0 0 7350 3850
use ddaa_slice  ddaa_slice_1
timestamp 1726841226
transform 1 0 7750 0 -1 11550
box 0 0 7350 3850
use ddaa_slice  ddaa_slice_2
timestamp 1726841226
transform 1 0 7750 0 1 11550
box 0 0 7350 3850
use ddaa_slice  ddaa_slice_3
timestamp 1726841226
transform 1 0 14950 0 1 11550
box 0 0 7350 3850
use ddaa_slice  ddaa_slice_4
timestamp 1726841226
transform 1 0 550 0 -1 11550
box 0 0 7350 3850
use ddaa_slice  ddaa_slice_5
timestamp 1726841226
transform 1 0 14950 0 -1 11550
box 0 0 7350 3850
use invdummy  invdummy_0
timestamp 1722856725
transform 1 0 22200 0 1 11550
box -50 0 300 3850
use invdummy  invdummy_1
timestamp 1722856725
transform -1 0 650 0 1 7700
box -50 0 300 3850
use invdummy  invdummy_5
timestamp 1722856725
transform -1 0 650 0 1 11550
box -50 0 300 3850
use invdummy  invdummy_6
timestamp 1722856725
transform 1 0 22200 0 1 7700
box -50 0 300 3850
use invedge  invedge_0
timestamp 1722865417
transform 1 0 22250 0 1 10450
box 150 1100 600 4950
use invedge  invedge_1
timestamp 1722865417
transform -1 0 600 0 1 6600
box 150 1100 600 4950
use invedge  invedge_5
timestamp 1722865417
transform -1 0 600 0 1 10450
box 150 1100 600 4950
use invedge  invedge_6
timestamp 1722865417
transform 1 0 22250 0 1 6600
box 150 1100 600 4950
<< labels >>
rlabel metal4 -800 15350 -750 15400 0 ipa
port 1 nsew
rlabel metal4 -600 15350 -550 15400 0 ima
port 2 nsew
rlabel metal4 -400 15350 -350 15400 0 ipb
port 3 nsew
rlabel metal4 -200 15350 -150 15400 0 imb
port 4 nsew
rlabel metal4 23400 15350 23650 15400 0 op
port 5 nsew
rlabel metal4 23000 15350 23250 15400 0 om
port 6 nsew
rlabel metal4 150 15350 200 15400 0 bp
port 7 nsew
rlabel metal4 300 15350 350 15400 0 bn
port 8 nsew
rlabel metal4 -1200 15350 -950 15400 0 vdd
port 9 nsew
rlabel metal4 -900 15350 -850 15400 0 vss
port 10 nsew
rlabel metal4 -1300 15350 -1250 15400 0 vsub
port 11 nsew
<< end >>
