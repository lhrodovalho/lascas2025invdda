magic
tech sky130A
timestamp 1726445033
<< locali >>
rect 50 3800 7300 3850
rect 50 2900 7300 2950
rect 50 2750 7300 2800
rect 50 1050 7300 1100
rect 50 900 7300 950
rect 50 0 7300 50
<< viali >>
rect 2765 2615 2785 2635
rect 4565 1215 4585 1235
rect 6365 1215 6385 1235
<< metal1 >>
rect 950 2640 1000 2650
rect 950 2610 960 2640
rect 990 2610 1000 2640
rect 950 2600 1000 2610
rect 2750 2640 2800 2650
rect 2750 2610 2760 2640
rect 2790 2610 2800 2640
rect 2750 2600 2800 2610
rect 4550 1240 4600 1250
rect 4550 1210 4560 1240
rect 4590 1210 4600 1240
rect 4550 1200 4600 1210
rect 6350 1240 6400 1250
rect 6350 1210 6360 1240
rect 6390 1210 6400 1240
rect 6350 1200 6400 1210
<< via1 >>
rect 960 2610 990 2640
rect 2760 2610 2790 2640
rect 4560 1235 4590 1240
rect 4560 1215 4565 1235
rect 4565 1215 4585 1235
rect 4585 1215 4590 1235
rect 4560 1210 4590 1215
rect 6360 1235 6390 1240
rect 6360 1215 6365 1235
rect 6365 1215 6385 1235
rect 6385 1215 6390 1235
rect 6360 1210 6390 1215
<< metal2 >>
rect 950 2640 1000 2650
rect 950 2610 960 2640
rect 990 2610 1000 2640
rect 950 2600 1000 2610
rect 2750 2640 2800 2650
rect 2750 2610 2760 2640
rect 2790 2610 2800 2640
rect 2750 2600 2800 2610
rect 4550 1240 4600 1250
rect 4550 1210 4560 1240
rect 4590 1210 4600 1240
rect 4550 1200 4600 1210
rect 6350 1240 6400 1250
rect 6350 1210 6360 1240
rect 6390 1210 6400 1240
rect 6350 1200 6400 1210
<< via2 >>
rect 960 2610 990 2640
rect 2760 2610 2790 2640
rect 4560 1210 4590 1240
rect 6360 1210 6390 1240
<< metal3 >>
rect 50 3700 7300 3750
rect 50 2800 7300 2850
rect 50 2700 7300 2750
rect 50 2645 7300 2650
rect 50 2640 2305 2645
rect 50 2610 960 2640
rect 990 2610 2305 2640
rect 50 2605 2305 2610
rect 2345 2640 5905 2645
rect 2345 2610 2760 2640
rect 2790 2610 5905 2640
rect 2345 2605 5905 2610
rect 5945 2605 7300 2645
rect 50 2600 7300 2605
rect 50 2500 7300 2550
rect 50 2300 7300 2350
rect 50 2145 7300 2150
rect 50 2105 505 2145
rect 545 2105 3205 2145
rect 3245 2105 7300 2145
rect 50 2100 7300 2105
rect 50 1745 7300 1750
rect 50 1705 4105 1745
rect 4145 1705 6805 1745
rect 6845 1705 7300 1745
rect 50 1700 7300 1705
rect 50 1300 7300 1350
rect 50 1245 7300 1250
rect 50 1205 1405 1245
rect 1445 1240 5005 1245
rect 1445 1210 4560 1240
rect 4590 1210 5005 1240
rect 1445 1205 5005 1210
rect 5045 1240 7300 1245
rect 5045 1210 6360 1240
rect 6390 1210 7300 1240
rect 5045 1205 7300 1210
rect 50 1200 7300 1205
rect 50 1100 7300 1150
rect 50 1000 7300 1050
rect 50 100 7300 150
<< via3 >>
rect 2305 2605 2345 2645
rect 5905 2605 5945 2645
rect 505 2105 545 2145
rect 3205 2105 3245 2145
rect 4105 1705 4145 1745
rect 6805 1705 6845 1745
rect 1405 1205 1445 1245
rect 5005 1205 5045 1245
<< metal4 >>
rect 2300 2645 2350 2650
rect 2300 2605 2305 2645
rect 2345 2605 2350 2645
rect 2300 2600 2350 2605
rect 5900 2645 5950 2650
rect 5900 2605 5905 2645
rect 5945 2605 5950 2645
rect 5900 2600 5950 2605
rect 500 2145 550 2150
rect 500 2105 505 2145
rect 545 2105 550 2145
rect 500 2100 550 2105
rect 3200 2145 3250 2150
rect 3200 2105 3205 2145
rect 3245 2105 3250 2145
rect 3200 2100 3250 2105
rect 4100 1745 4150 1750
rect 4100 1705 4105 1745
rect 4145 1705 4150 1745
rect 4100 1700 4150 1705
rect 6800 1745 6850 1750
rect 6800 1705 6805 1745
rect 6845 1705 6850 1745
rect 6800 1700 6850 1705
rect 1400 1245 1450 1250
rect 1400 1205 1405 1245
rect 1445 1205 1450 1245
rect 1400 1200 1450 1205
rect 5000 1245 5050 1250
rect 5000 1205 5005 1245
rect 5045 1205 5050 1245
rect 5000 1200 5050 1205
use inv1p1  a0
timestamp 1726000395
transform 1 0 50 0 1 0
box -50 0 1000 3850
use inv1p1  a1
timestamp 1726000395
transform -1 0 1900 0 1 0
box -50 0 1000 3850
use inv1p1  a2
timestamp 1726000395
transform 1 0 1850 0 1 0
box -50 0 1000 3850
use inv1p1  a3
timestamp 1726000395
transform -1 0 3700 0 1 0
box -50 0 1000 3850
use inv1p1  a4
timestamp 1726000395
transform 1 0 3650 0 1 0
box -50 0 1000 3850
use inv1p1  a5
timestamp 1726000395
transform -1 0 5500 0 1 0
box -50 0 1000 3850
use inv1p1  a6
timestamp 1726000395
transform 1 0 5450 0 1 0
box -50 0 1000 3850
use inv1p1  a7
timestamp 1726000395
transform -1 0 7300 0 1 0
box -50 0 1000 3850
<< labels >>
rlabel metal3 50 2100 7300 2150 0 ip
port 1 nsew
rlabel metal3 50 1700 7300 1750 0 im
port 2 nsew
rlabel metal3 50 2600 7300 2650 0 xm
port 3 nsew
rlabel metal3 50 1200 7300 1250 0 xp
port 4 nsew
rlabel metal3 50 2700 7300 2750 0 op
port 5 nsew
rlabel metal3 50 2500 7300 2550 0 op
port 5 nsew
rlabel metal3 50 1300 7300 1350 0 om
port 6 nsew
rlabel metal3 50 1100 7300 1150 0 om
port 6 nsew
rlabel locali 50 2900 7300 2950 0 bp
port 7 nsew
rlabel locali 50 900 7300 950 0 bp
port 7 nsew
rlabel locali 50 2750 7300 2800 0 bn
port 8 nsew
rlabel locali 50 1050 7300 1100 0 bn
port 8 nsew
rlabel metal3 50 3700 7300 3750 0 vdd
port 9 nsew
rlabel metal3 50 100 7300 150 0 vdd
port 9 nsew
rlabel metal3 50 2800 7300 2850 0 vss
port 10 nsew
rlabel metal3 50 1000 7300 1050 0 vss
port 10 nsew
rlabel locali 50 3800 7300 3850 0 vsub
port 11 nsew
rlabel locali 50 0 7300 50 0 vsub
port 11 nsew
<< end >>
