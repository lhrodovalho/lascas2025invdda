magic
tech sky130A
timestamp 1726000395
<< dnwell >>
rect 0 895 950 2955
<< nwell >>
rect -50 2850 1000 3750
rect -50 100 1000 1000
<< pwell >>
rect 0 2000 950 2850
rect 0 1850 900 2000
rect 0 1000 950 1850
<< nmos >>
rect 50 2000 450 2700
rect 500 2000 900 2700
rect 50 1150 450 1850
rect 500 1150 900 1850
<< pmoslvt >>
rect 50 3100 450 3600
rect 500 3100 900 3600
rect 50 250 450 750
rect 500 250 900 750
<< ndiff >>
rect 0 2685 50 2700
rect 0 2665 15 2685
rect 35 2665 50 2685
rect 0 2635 50 2665
rect 0 2615 15 2635
rect 35 2615 50 2635
rect 0 2585 50 2615
rect 0 2565 15 2585
rect 35 2565 50 2585
rect 0 2535 50 2565
rect 0 2515 15 2535
rect 35 2515 50 2535
rect 0 2485 50 2515
rect 0 2465 15 2485
rect 35 2465 50 2485
rect 0 2435 50 2465
rect 0 2415 15 2435
rect 35 2415 50 2435
rect 0 2385 50 2415
rect 0 2365 15 2385
rect 35 2365 50 2385
rect 0 2335 50 2365
rect 0 2315 15 2335
rect 35 2315 50 2335
rect 0 2285 50 2315
rect 0 2265 15 2285
rect 35 2265 50 2285
rect 0 2235 50 2265
rect 0 2215 15 2235
rect 35 2215 50 2235
rect 0 2185 50 2215
rect 0 2165 15 2185
rect 35 2165 50 2185
rect 0 2135 50 2165
rect 0 2115 15 2135
rect 35 2115 50 2135
rect 0 2085 50 2115
rect 0 2065 15 2085
rect 35 2065 50 2085
rect 0 2035 50 2065
rect 0 2015 15 2035
rect 35 2015 50 2035
rect 0 2000 50 2015
rect 450 2000 500 2700
rect 900 2685 950 2700
rect 900 2665 915 2685
rect 935 2665 950 2685
rect 900 2635 950 2665
rect 900 2615 915 2635
rect 935 2615 950 2635
rect 900 2585 950 2615
rect 900 2565 915 2585
rect 935 2565 950 2585
rect 900 2535 950 2565
rect 900 2515 915 2535
rect 935 2515 950 2535
rect 900 2485 950 2515
rect 900 2465 915 2485
rect 935 2465 950 2485
rect 900 2435 950 2465
rect 900 2415 915 2435
rect 935 2415 950 2435
rect 900 2385 950 2415
rect 900 2365 915 2385
rect 935 2365 950 2385
rect 900 2335 950 2365
rect 900 2315 915 2335
rect 935 2315 950 2335
rect 900 2285 950 2315
rect 900 2265 915 2285
rect 935 2265 950 2285
rect 900 2235 950 2265
rect 900 2215 915 2235
rect 935 2215 950 2235
rect 900 2185 950 2215
rect 900 2165 915 2185
rect 935 2165 950 2185
rect 900 2135 950 2165
rect 900 2115 915 2135
rect 935 2115 950 2135
rect 900 2085 950 2115
rect 900 2065 915 2085
rect 935 2065 950 2085
rect 900 2035 950 2065
rect 900 2015 915 2035
rect 935 2015 950 2035
rect 900 2000 950 2015
rect 0 1835 50 1850
rect 0 1815 15 1835
rect 35 1815 50 1835
rect 0 1785 50 1815
rect 0 1765 15 1785
rect 35 1765 50 1785
rect 0 1735 50 1765
rect 0 1715 15 1735
rect 35 1715 50 1735
rect 0 1685 50 1715
rect 0 1665 15 1685
rect 35 1665 50 1685
rect 0 1635 50 1665
rect 0 1615 15 1635
rect 35 1615 50 1635
rect 0 1585 50 1615
rect 0 1565 15 1585
rect 35 1565 50 1585
rect 0 1535 50 1565
rect 0 1515 15 1535
rect 35 1515 50 1535
rect 0 1485 50 1515
rect 0 1465 15 1485
rect 35 1465 50 1485
rect 0 1435 50 1465
rect 0 1415 15 1435
rect 35 1415 50 1435
rect 0 1385 50 1415
rect 0 1365 15 1385
rect 35 1365 50 1385
rect 0 1335 50 1365
rect 0 1315 15 1335
rect 35 1315 50 1335
rect 0 1285 50 1315
rect 0 1265 15 1285
rect 35 1265 50 1285
rect 0 1235 50 1265
rect 0 1215 15 1235
rect 35 1215 50 1235
rect 0 1185 50 1215
rect 0 1165 15 1185
rect 35 1165 50 1185
rect 0 1150 50 1165
rect 450 1150 500 1850
rect 900 1835 950 1850
rect 900 1815 915 1835
rect 935 1815 950 1835
rect 900 1785 950 1815
rect 900 1765 915 1785
rect 935 1765 950 1785
rect 900 1735 950 1765
rect 900 1715 915 1735
rect 935 1715 950 1735
rect 900 1685 950 1715
rect 900 1665 915 1685
rect 935 1665 950 1685
rect 900 1635 950 1665
rect 900 1615 915 1635
rect 935 1615 950 1635
rect 900 1585 950 1615
rect 900 1565 915 1585
rect 935 1565 950 1585
rect 900 1535 950 1565
rect 900 1515 915 1535
rect 935 1515 950 1535
rect 900 1485 950 1515
rect 900 1465 915 1485
rect 935 1465 950 1485
rect 900 1435 950 1465
rect 900 1415 915 1435
rect 935 1415 950 1435
rect 900 1385 950 1415
rect 900 1365 915 1385
rect 935 1365 950 1385
rect 900 1335 950 1365
rect 900 1315 915 1335
rect 935 1315 950 1335
rect 900 1285 950 1315
rect 900 1265 915 1285
rect 935 1265 950 1285
rect 900 1235 950 1265
rect 900 1215 915 1235
rect 935 1215 950 1235
rect 900 1185 950 1215
rect 900 1165 915 1185
rect 935 1165 950 1185
rect 900 1150 950 1165
<< pdiff >>
rect 0 3585 50 3600
rect 0 3565 15 3585
rect 35 3565 50 3585
rect 0 3535 50 3565
rect 0 3515 15 3535
rect 35 3515 50 3535
rect 0 3485 50 3515
rect 0 3465 15 3485
rect 35 3465 50 3485
rect 0 3435 50 3465
rect 0 3415 15 3435
rect 35 3415 50 3435
rect 0 3385 50 3415
rect 0 3365 15 3385
rect 35 3365 50 3385
rect 0 3335 50 3365
rect 0 3315 15 3335
rect 35 3315 50 3335
rect 0 3285 50 3315
rect 0 3265 15 3285
rect 35 3265 50 3285
rect 0 3235 50 3265
rect 0 3215 15 3235
rect 35 3215 50 3235
rect 0 3185 50 3215
rect 0 3165 15 3185
rect 35 3165 50 3185
rect 0 3135 50 3165
rect 0 3115 15 3135
rect 35 3115 50 3135
rect 0 3100 50 3115
rect 450 3585 500 3600
rect 450 3565 465 3585
rect 485 3565 500 3585
rect 450 3535 500 3565
rect 450 3515 465 3535
rect 485 3515 500 3535
rect 450 3485 500 3515
rect 450 3465 465 3485
rect 485 3465 500 3485
rect 450 3435 500 3465
rect 450 3415 465 3435
rect 485 3415 500 3435
rect 450 3385 500 3415
rect 450 3365 465 3385
rect 485 3365 500 3385
rect 450 3335 500 3365
rect 450 3315 465 3335
rect 485 3315 500 3335
rect 450 3285 500 3315
rect 450 3265 465 3285
rect 485 3265 500 3285
rect 450 3235 500 3265
rect 450 3215 465 3235
rect 485 3215 500 3235
rect 450 3185 500 3215
rect 450 3165 465 3185
rect 485 3165 500 3185
rect 450 3135 500 3165
rect 450 3115 465 3135
rect 485 3115 500 3135
rect 450 3100 500 3115
rect 900 3585 950 3600
rect 900 3565 915 3585
rect 935 3565 950 3585
rect 900 3535 950 3565
rect 900 3515 915 3535
rect 935 3515 950 3535
rect 900 3485 950 3515
rect 900 3465 915 3485
rect 935 3465 950 3485
rect 900 3435 950 3465
rect 900 3415 915 3435
rect 935 3415 950 3435
rect 900 3385 950 3415
rect 900 3365 915 3385
rect 935 3365 950 3385
rect 900 3335 950 3365
rect 900 3315 915 3335
rect 935 3315 950 3335
rect 900 3285 950 3315
rect 900 3265 915 3285
rect 935 3265 950 3285
rect 900 3235 950 3265
rect 900 3215 915 3235
rect 935 3215 950 3235
rect 900 3185 950 3215
rect 900 3165 915 3185
rect 935 3165 950 3185
rect 900 3135 950 3165
rect 900 3115 915 3135
rect 935 3115 950 3135
rect 900 3100 950 3115
rect 0 735 50 750
rect 0 715 15 735
rect 35 715 50 735
rect 0 685 50 715
rect 0 665 15 685
rect 35 665 50 685
rect 0 635 50 665
rect 0 615 15 635
rect 35 615 50 635
rect 0 585 50 615
rect 0 565 15 585
rect 35 565 50 585
rect 0 535 50 565
rect 0 515 15 535
rect 35 515 50 535
rect 0 485 50 515
rect 0 465 15 485
rect 35 465 50 485
rect 0 435 50 465
rect 0 415 15 435
rect 35 415 50 435
rect 0 385 50 415
rect 0 365 15 385
rect 35 365 50 385
rect 0 335 50 365
rect 0 315 15 335
rect 35 315 50 335
rect 0 285 50 315
rect 0 265 15 285
rect 35 265 50 285
rect 0 250 50 265
rect 450 735 500 750
rect 450 715 465 735
rect 485 715 500 735
rect 450 685 500 715
rect 450 665 465 685
rect 485 665 500 685
rect 450 635 500 665
rect 450 615 465 635
rect 485 615 500 635
rect 450 585 500 615
rect 450 565 465 585
rect 485 565 500 585
rect 450 535 500 565
rect 450 515 465 535
rect 485 515 500 535
rect 450 485 500 515
rect 450 465 465 485
rect 485 465 500 485
rect 450 435 500 465
rect 450 415 465 435
rect 485 415 500 435
rect 450 385 500 415
rect 450 365 465 385
rect 485 365 500 385
rect 450 335 500 365
rect 450 315 465 335
rect 485 315 500 335
rect 450 285 500 315
rect 450 265 465 285
rect 485 265 500 285
rect 450 250 500 265
rect 900 735 950 750
rect 900 715 915 735
rect 935 715 950 735
rect 900 685 950 715
rect 900 665 915 685
rect 935 665 950 685
rect 900 635 950 665
rect 900 615 915 635
rect 935 615 950 635
rect 900 585 950 615
rect 900 565 915 585
rect 935 565 950 585
rect 900 535 950 565
rect 900 515 915 535
rect 935 515 950 535
rect 900 485 950 515
rect 900 465 915 485
rect 935 465 950 485
rect 900 435 950 465
rect 900 415 915 435
rect 935 415 950 435
rect 900 385 950 415
rect 900 365 915 385
rect 935 365 950 385
rect 900 335 950 365
rect 900 315 915 335
rect 935 315 950 335
rect 900 285 950 315
rect 900 265 915 285
rect 935 265 950 285
rect 900 250 950 265
<< ndiffc >>
rect 15 2665 35 2685
rect 15 2615 35 2635
rect 15 2565 35 2585
rect 15 2515 35 2535
rect 15 2465 35 2485
rect 15 2415 35 2435
rect 15 2365 35 2385
rect 15 2315 35 2335
rect 15 2265 35 2285
rect 15 2215 35 2235
rect 15 2165 35 2185
rect 15 2115 35 2135
rect 15 2065 35 2085
rect 15 2015 35 2035
rect 915 2665 935 2685
rect 915 2615 935 2635
rect 915 2565 935 2585
rect 915 2515 935 2535
rect 915 2465 935 2485
rect 915 2415 935 2435
rect 915 2365 935 2385
rect 915 2315 935 2335
rect 915 2265 935 2285
rect 915 2215 935 2235
rect 915 2165 935 2185
rect 915 2115 935 2135
rect 915 2065 935 2085
rect 915 2015 935 2035
rect 15 1815 35 1835
rect 15 1765 35 1785
rect 15 1715 35 1735
rect 15 1665 35 1685
rect 15 1615 35 1635
rect 15 1565 35 1585
rect 15 1515 35 1535
rect 15 1465 35 1485
rect 15 1415 35 1435
rect 15 1365 35 1385
rect 15 1315 35 1335
rect 15 1265 35 1285
rect 15 1215 35 1235
rect 15 1165 35 1185
rect 915 1815 935 1835
rect 915 1765 935 1785
rect 915 1715 935 1735
rect 915 1665 935 1685
rect 915 1615 935 1635
rect 915 1565 935 1585
rect 915 1515 935 1535
rect 915 1465 935 1485
rect 915 1415 935 1435
rect 915 1365 935 1385
rect 915 1315 935 1335
rect 915 1265 935 1285
rect 915 1215 935 1235
rect 915 1165 935 1185
<< pdiffc >>
rect 15 3565 35 3585
rect 15 3515 35 3535
rect 15 3465 35 3485
rect 15 3415 35 3435
rect 15 3365 35 3385
rect 15 3315 35 3335
rect 15 3265 35 3285
rect 15 3215 35 3235
rect 15 3165 35 3185
rect 15 3115 35 3135
rect 465 3565 485 3585
rect 465 3515 485 3535
rect 465 3465 485 3485
rect 465 3415 485 3435
rect 465 3365 485 3385
rect 465 3315 485 3335
rect 465 3265 485 3285
rect 465 3215 485 3235
rect 465 3165 485 3185
rect 465 3115 485 3135
rect 915 3565 935 3585
rect 915 3515 935 3535
rect 915 3465 935 3485
rect 915 3415 935 3435
rect 915 3365 935 3385
rect 915 3315 935 3335
rect 915 3265 935 3285
rect 915 3215 935 3235
rect 915 3165 935 3185
rect 915 3115 935 3135
rect 15 715 35 735
rect 15 665 35 685
rect 15 615 35 635
rect 15 565 35 585
rect 15 515 35 535
rect 15 465 35 485
rect 15 415 35 435
rect 15 365 35 385
rect 15 315 35 335
rect 15 265 35 285
rect 465 715 485 735
rect 465 665 485 685
rect 465 615 485 635
rect 465 565 485 585
rect 465 515 485 535
rect 465 465 485 485
rect 465 415 485 435
rect 465 365 485 385
rect 465 315 485 335
rect 465 265 485 285
rect 915 715 935 735
rect 915 665 935 685
rect 915 615 935 635
rect 915 565 935 585
rect 915 515 935 535
rect 915 465 935 485
rect 915 415 935 435
rect 915 365 935 385
rect 915 315 935 335
rect 915 265 935 285
<< psubdiff >>
rect 0 3835 950 3850
rect 0 3815 15 3835
rect 35 3815 65 3835
rect 85 3815 115 3835
rect 135 3815 165 3835
rect 185 3815 215 3835
rect 235 3815 265 3835
rect 285 3815 315 3835
rect 335 3815 365 3835
rect 385 3815 415 3835
rect 435 3815 465 3835
rect 485 3815 515 3835
rect 535 3815 565 3835
rect 585 3815 615 3835
rect 635 3815 665 3835
rect 685 3815 715 3835
rect 735 3815 765 3835
rect 785 3815 815 3835
rect 835 3815 865 3835
rect 885 3815 915 3835
rect 935 3815 950 3835
rect 0 3800 950 3815
rect 0 2785 950 2800
rect 0 2765 15 2785
rect 35 2765 65 2785
rect 85 2765 115 2785
rect 135 2765 165 2785
rect 185 2765 215 2785
rect 235 2765 265 2785
rect 285 2765 315 2785
rect 335 2765 365 2785
rect 385 2765 415 2785
rect 435 2765 465 2785
rect 485 2765 515 2785
rect 535 2765 565 2785
rect 585 2765 615 2785
rect 635 2765 665 2785
rect 685 2765 715 2785
rect 735 2765 765 2785
rect 785 2765 815 2785
rect 835 2765 865 2785
rect 885 2765 915 2785
rect 935 2765 950 2785
rect 0 2750 950 2765
rect 0 1085 950 1100
rect 0 1065 15 1085
rect 35 1065 65 1085
rect 85 1065 115 1085
rect 135 1065 165 1085
rect 185 1065 215 1085
rect 235 1065 265 1085
rect 285 1065 315 1085
rect 335 1065 365 1085
rect 385 1065 415 1085
rect 435 1065 465 1085
rect 485 1065 515 1085
rect 535 1065 565 1085
rect 585 1065 615 1085
rect 635 1065 665 1085
rect 685 1065 715 1085
rect 735 1065 765 1085
rect 785 1065 815 1085
rect 835 1065 865 1085
rect 885 1065 915 1085
rect 935 1065 950 1085
rect 0 1050 950 1065
rect 0 35 950 50
rect 0 15 15 35
rect 35 15 65 35
rect 85 15 115 35
rect 135 15 165 35
rect 185 15 215 35
rect 235 15 265 35
rect 285 15 315 35
rect 335 15 365 35
rect 385 15 415 35
rect 435 15 465 35
rect 485 15 515 35
rect 535 15 565 35
rect 585 15 615 35
rect 635 15 665 35
rect 685 15 715 35
rect 735 15 765 35
rect 785 15 815 35
rect 835 15 865 35
rect 885 15 915 35
rect 935 15 950 35
rect 0 0 950 15
<< nsubdiff >>
rect 0 3685 950 3700
rect 0 3665 15 3685
rect 35 3665 65 3685
rect 85 3665 115 3685
rect 135 3665 165 3685
rect 185 3665 215 3685
rect 235 3665 265 3685
rect 285 3665 315 3685
rect 335 3665 365 3685
rect 385 3665 415 3685
rect 435 3665 465 3685
rect 485 3665 515 3685
rect 535 3665 565 3685
rect 585 3665 615 3685
rect 635 3665 665 3685
rect 685 3665 715 3685
rect 735 3665 765 3685
rect 785 3665 815 3685
rect 835 3665 865 3685
rect 885 3665 915 3685
rect 935 3665 950 3685
rect 0 3650 950 3665
rect 0 2935 950 2950
rect 0 2915 15 2935
rect 35 2915 65 2935
rect 85 2915 115 2935
rect 135 2915 165 2935
rect 185 2915 215 2935
rect 235 2915 265 2935
rect 285 2915 315 2935
rect 335 2915 365 2935
rect 385 2915 415 2935
rect 435 2915 465 2935
rect 485 2915 515 2935
rect 535 2915 565 2935
rect 585 2915 615 2935
rect 635 2915 665 2935
rect 685 2915 715 2935
rect 735 2915 765 2935
rect 785 2915 815 2935
rect 835 2915 865 2935
rect 885 2915 915 2935
rect 935 2915 950 2935
rect 0 2900 950 2915
rect 0 935 950 950
rect 0 915 15 935
rect 35 915 65 935
rect 85 915 115 935
rect 135 915 165 935
rect 185 915 215 935
rect 235 915 265 935
rect 285 915 315 935
rect 335 915 365 935
rect 385 915 415 935
rect 435 915 465 935
rect 485 915 515 935
rect 535 915 565 935
rect 585 915 615 935
rect 635 915 665 935
rect 685 915 715 935
rect 735 915 765 935
rect 785 915 815 935
rect 835 915 865 935
rect 885 915 915 935
rect 935 915 950 935
rect 0 900 950 915
rect 0 185 950 200
rect 0 165 15 185
rect 35 165 65 185
rect 85 165 115 185
rect 135 165 165 185
rect 185 165 215 185
rect 235 165 265 185
rect 285 165 315 185
rect 335 165 365 185
rect 385 165 415 185
rect 435 165 465 185
rect 485 165 515 185
rect 535 165 565 185
rect 585 165 615 185
rect 635 165 665 185
rect 685 165 715 185
rect 735 165 765 185
rect 785 165 815 185
rect 835 165 865 185
rect 885 165 915 185
rect 935 165 950 185
rect 0 150 950 165
<< psubdiffcont >>
rect 15 3815 35 3835
rect 65 3815 85 3835
rect 115 3815 135 3835
rect 165 3815 185 3835
rect 215 3815 235 3835
rect 265 3815 285 3835
rect 315 3815 335 3835
rect 365 3815 385 3835
rect 415 3815 435 3835
rect 465 3815 485 3835
rect 515 3815 535 3835
rect 565 3815 585 3835
rect 615 3815 635 3835
rect 665 3815 685 3835
rect 715 3815 735 3835
rect 765 3815 785 3835
rect 815 3815 835 3835
rect 865 3815 885 3835
rect 915 3815 935 3835
rect 15 2765 35 2785
rect 65 2765 85 2785
rect 115 2765 135 2785
rect 165 2765 185 2785
rect 215 2765 235 2785
rect 265 2765 285 2785
rect 315 2765 335 2785
rect 365 2765 385 2785
rect 415 2765 435 2785
rect 465 2765 485 2785
rect 515 2765 535 2785
rect 565 2765 585 2785
rect 615 2765 635 2785
rect 665 2765 685 2785
rect 715 2765 735 2785
rect 765 2765 785 2785
rect 815 2765 835 2785
rect 865 2765 885 2785
rect 915 2765 935 2785
rect 15 1065 35 1085
rect 65 1065 85 1085
rect 115 1065 135 1085
rect 165 1065 185 1085
rect 215 1065 235 1085
rect 265 1065 285 1085
rect 315 1065 335 1085
rect 365 1065 385 1085
rect 415 1065 435 1085
rect 465 1065 485 1085
rect 515 1065 535 1085
rect 565 1065 585 1085
rect 615 1065 635 1085
rect 665 1065 685 1085
rect 715 1065 735 1085
rect 765 1065 785 1085
rect 815 1065 835 1085
rect 865 1065 885 1085
rect 915 1065 935 1085
rect 15 15 35 35
rect 65 15 85 35
rect 115 15 135 35
rect 165 15 185 35
rect 215 15 235 35
rect 265 15 285 35
rect 315 15 335 35
rect 365 15 385 35
rect 415 15 435 35
rect 465 15 485 35
rect 515 15 535 35
rect 565 15 585 35
rect 615 15 635 35
rect 665 15 685 35
rect 715 15 735 35
rect 765 15 785 35
rect 815 15 835 35
rect 865 15 885 35
rect 915 15 935 35
<< nsubdiffcont >>
rect 15 3665 35 3685
rect 65 3665 85 3685
rect 115 3665 135 3685
rect 165 3665 185 3685
rect 215 3665 235 3685
rect 265 3665 285 3685
rect 315 3665 335 3685
rect 365 3665 385 3685
rect 415 3665 435 3685
rect 465 3665 485 3685
rect 515 3665 535 3685
rect 565 3665 585 3685
rect 615 3665 635 3685
rect 665 3665 685 3685
rect 715 3665 735 3685
rect 765 3665 785 3685
rect 815 3665 835 3685
rect 865 3665 885 3685
rect 915 3665 935 3685
rect 15 2915 35 2935
rect 65 2915 85 2935
rect 115 2915 135 2935
rect 165 2915 185 2935
rect 215 2915 235 2935
rect 265 2915 285 2935
rect 315 2915 335 2935
rect 365 2915 385 2935
rect 415 2915 435 2935
rect 465 2915 485 2935
rect 515 2915 535 2935
rect 565 2915 585 2935
rect 615 2915 635 2935
rect 665 2915 685 2935
rect 715 2915 735 2935
rect 765 2915 785 2935
rect 815 2915 835 2935
rect 865 2915 885 2935
rect 915 2915 935 2935
rect 15 915 35 935
rect 65 915 85 935
rect 115 915 135 935
rect 165 915 185 935
rect 215 915 235 935
rect 265 915 285 935
rect 315 915 335 935
rect 365 915 385 935
rect 415 915 435 935
rect 465 915 485 935
rect 515 915 535 935
rect 565 915 585 935
rect 615 915 635 935
rect 665 915 685 935
rect 715 915 735 935
rect 765 915 785 935
rect 815 915 835 935
rect 865 915 885 935
rect 915 915 935 935
rect 15 165 35 185
rect 65 165 85 185
rect 115 165 135 185
rect 165 165 185 185
rect 215 165 235 185
rect 265 165 285 185
rect 315 165 335 185
rect 365 165 385 185
rect 415 165 435 185
rect 465 165 485 185
rect 515 165 535 185
rect 565 165 585 185
rect 615 165 635 185
rect 665 165 685 185
rect 715 165 735 185
rect 765 165 785 185
rect 815 165 835 185
rect 865 165 885 185
rect 915 165 935 185
<< poly >>
rect 50 3600 450 3615
rect 500 3600 900 3615
rect 50 3050 450 3100
rect 500 3050 900 3100
rect 50 3035 900 3050
rect 50 3015 65 3035
rect 85 3015 115 3035
rect 135 3015 165 3035
rect 185 3015 215 3035
rect 235 3015 265 3035
rect 285 3015 315 3035
rect 335 3015 365 3035
rect 385 3015 415 3035
rect 435 3015 465 3035
rect 485 3015 515 3035
rect 535 3015 565 3035
rect 585 3015 615 3035
rect 635 3015 665 3035
rect 685 3015 715 3035
rect 735 3015 765 3035
rect 785 3015 815 3035
rect 835 3015 865 3035
rect 885 3015 900 3035
rect 50 3000 900 3015
rect 50 2700 450 2715
rect 500 2700 900 2715
rect 50 1950 450 2000
rect 500 1950 900 2000
rect 50 1935 900 1950
rect 50 1915 65 1935
rect 85 1915 115 1935
rect 135 1915 165 1935
rect 185 1915 215 1935
rect 235 1915 265 1935
rect 285 1915 315 1935
rect 335 1915 365 1935
rect 385 1915 415 1935
rect 435 1915 465 1935
rect 485 1915 515 1935
rect 535 1915 565 1935
rect 585 1915 615 1935
rect 635 1915 665 1935
rect 685 1915 715 1935
rect 735 1915 765 1935
rect 785 1915 815 1935
rect 835 1915 865 1935
rect 885 1915 900 1935
rect 50 1900 900 1915
rect 50 1850 450 1900
rect 500 1850 900 1900
rect 50 1135 450 1150
rect 500 1135 900 1150
rect 50 835 900 850
rect 50 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 215 835
rect 235 815 265 835
rect 285 815 315 835
rect 335 815 365 835
rect 385 815 415 835
rect 435 815 465 835
rect 485 815 515 835
rect 535 815 565 835
rect 585 815 615 835
rect 635 815 665 835
rect 685 815 715 835
rect 735 815 765 835
rect 785 815 815 835
rect 835 815 865 835
rect 885 815 900 835
rect 50 800 900 815
rect 50 750 450 800
rect 500 750 900 800
rect 50 235 450 250
rect 500 235 900 250
<< polycont >>
rect 65 3015 85 3035
rect 115 3015 135 3035
rect 165 3015 185 3035
rect 215 3015 235 3035
rect 265 3015 285 3035
rect 315 3015 335 3035
rect 365 3015 385 3035
rect 415 3015 435 3035
rect 465 3015 485 3035
rect 515 3015 535 3035
rect 565 3015 585 3035
rect 615 3015 635 3035
rect 665 3015 685 3035
rect 715 3015 735 3035
rect 765 3015 785 3035
rect 815 3015 835 3035
rect 865 3015 885 3035
rect 65 1915 85 1935
rect 115 1915 135 1935
rect 165 1915 185 1935
rect 215 1915 235 1935
rect 265 1915 285 1935
rect 315 1915 335 1935
rect 365 1915 385 1935
rect 415 1915 435 1935
rect 465 1915 485 1935
rect 515 1915 535 1935
rect 565 1915 585 1935
rect 615 1915 635 1935
rect 665 1915 685 1935
rect 715 1915 735 1935
rect 765 1915 785 1935
rect 815 1915 835 1935
rect 865 1915 885 1935
rect 65 815 85 835
rect 115 815 135 835
rect 165 815 185 835
rect 215 815 235 835
rect 265 815 285 835
rect 315 815 335 835
rect 365 815 385 835
rect 415 815 435 835
rect 465 815 485 835
rect 515 815 535 835
rect 565 815 585 835
rect 615 815 635 835
rect 665 815 685 835
rect 715 815 735 835
rect 765 815 785 835
rect 815 815 835 835
rect 865 815 885 835
<< locali >>
rect 0 3835 950 3850
rect 0 3815 15 3835
rect 35 3815 65 3835
rect 85 3815 115 3835
rect 135 3815 165 3835
rect 185 3815 215 3835
rect 235 3815 265 3835
rect 285 3815 315 3835
rect 335 3815 365 3835
rect 385 3815 415 3835
rect 435 3815 465 3835
rect 485 3815 515 3835
rect 535 3815 565 3835
rect 585 3815 615 3835
rect 635 3815 665 3835
rect 685 3815 715 3835
rect 735 3815 765 3835
rect 785 3815 815 3835
rect 835 3815 865 3835
rect 885 3815 915 3835
rect 935 3815 950 3835
rect 0 3800 950 3815
rect 0 3685 950 3700
rect 0 3665 15 3685
rect 35 3665 65 3685
rect 85 3665 115 3685
rect 135 3665 165 3685
rect 185 3665 215 3685
rect 235 3665 265 3685
rect 285 3665 315 3685
rect 335 3665 365 3685
rect 385 3665 415 3685
rect 435 3665 465 3685
rect 485 3665 515 3685
rect 535 3665 565 3685
rect 585 3665 615 3685
rect 635 3665 665 3685
rect 685 3665 715 3685
rect 735 3665 765 3685
rect 785 3665 815 3685
rect 835 3665 865 3685
rect 885 3665 915 3685
rect 935 3665 950 3685
rect 0 3650 950 3665
rect 0 3585 50 3600
rect 0 3565 15 3585
rect 35 3565 50 3585
rect 0 3535 50 3565
rect 0 3515 15 3535
rect 35 3515 50 3535
rect 0 3485 50 3515
rect 0 3465 15 3485
rect 35 3465 50 3485
rect 0 3435 50 3465
rect 0 3415 15 3435
rect 35 3415 50 3435
rect 0 3385 50 3415
rect 0 3365 15 3385
rect 35 3365 50 3385
rect 0 3335 50 3365
rect 0 3315 15 3335
rect 35 3315 50 3335
rect 0 3285 50 3315
rect 0 3265 15 3285
rect 35 3265 50 3285
rect 0 3235 50 3265
rect 0 3215 15 3235
rect 35 3215 50 3235
rect 0 3185 50 3215
rect 0 3165 15 3185
rect 35 3165 50 3185
rect 0 3135 50 3165
rect 0 3115 15 3135
rect 35 3115 50 3135
rect 0 3100 50 3115
rect 450 3585 500 3600
rect 450 3565 465 3585
rect 485 3565 500 3585
rect 450 3535 500 3565
rect 450 3515 465 3535
rect 485 3515 500 3535
rect 450 3485 500 3515
rect 450 3465 465 3485
rect 485 3465 500 3485
rect 450 3435 500 3465
rect 450 3415 465 3435
rect 485 3415 500 3435
rect 450 3385 500 3415
rect 450 3365 465 3385
rect 485 3365 500 3385
rect 450 3335 500 3365
rect 450 3315 465 3335
rect 485 3315 500 3335
rect 450 3285 500 3315
rect 450 3265 465 3285
rect 485 3265 500 3285
rect 450 3235 500 3265
rect 450 3215 465 3235
rect 485 3215 500 3235
rect 450 3185 500 3215
rect 450 3165 465 3185
rect 485 3165 500 3185
rect 450 3135 500 3165
rect 450 3115 465 3135
rect 485 3115 500 3135
rect 450 3100 500 3115
rect 900 3585 950 3600
rect 900 3565 915 3585
rect 935 3565 950 3585
rect 900 3535 950 3565
rect 900 3515 915 3535
rect 935 3515 950 3535
rect 900 3485 950 3515
rect 900 3465 915 3485
rect 935 3465 950 3485
rect 900 3435 950 3465
rect 900 3415 915 3435
rect 935 3415 950 3435
rect 900 3385 950 3415
rect 900 3365 915 3385
rect 935 3365 950 3385
rect 900 3335 950 3365
rect 900 3315 915 3335
rect 935 3315 950 3335
rect 900 3285 950 3315
rect 900 3265 915 3285
rect 935 3265 950 3285
rect 900 3235 950 3265
rect 900 3215 915 3235
rect 935 3215 950 3235
rect 900 3185 950 3215
rect 900 3165 915 3185
rect 935 3165 950 3185
rect 900 3135 950 3165
rect 900 3115 915 3135
rect 935 3115 950 3135
rect 900 3100 950 3115
rect 50 3035 900 3050
rect 50 3015 65 3035
rect 85 3015 115 3035
rect 135 3015 165 3035
rect 185 3015 215 3035
rect 235 3015 265 3035
rect 285 3015 315 3035
rect 335 3015 365 3035
rect 385 3015 415 3035
rect 435 3015 465 3035
rect 485 3015 515 3035
rect 535 3015 565 3035
rect 585 3015 615 3035
rect 635 3015 665 3035
rect 685 3015 715 3035
rect 735 3015 765 3035
rect 785 3015 815 3035
rect 835 3015 865 3035
rect 885 3015 900 3035
rect 50 3000 900 3015
rect 0 2935 950 2950
rect 0 2915 15 2935
rect 35 2915 65 2935
rect 85 2915 115 2935
rect 135 2915 165 2935
rect 185 2915 215 2935
rect 235 2915 265 2935
rect 285 2915 315 2935
rect 335 2915 365 2935
rect 385 2915 415 2935
rect 435 2915 465 2935
rect 485 2915 515 2935
rect 535 2915 565 2935
rect 585 2915 615 2935
rect 635 2915 665 2935
rect 685 2915 715 2935
rect 735 2915 765 2935
rect 785 2915 815 2935
rect 835 2915 865 2935
rect 885 2915 915 2935
rect 935 2915 950 2935
rect 0 2900 950 2915
rect 0 2785 950 2800
rect 0 2765 15 2785
rect 35 2765 65 2785
rect 85 2765 115 2785
rect 135 2765 165 2785
rect 185 2765 215 2785
rect 235 2765 265 2785
rect 285 2765 315 2785
rect 335 2765 365 2785
rect 385 2765 415 2785
rect 435 2765 465 2785
rect 485 2765 515 2785
rect 535 2765 565 2785
rect 585 2765 615 2785
rect 635 2765 665 2785
rect 685 2765 715 2785
rect 735 2765 765 2785
rect 785 2765 815 2785
rect 835 2765 865 2785
rect 885 2765 915 2785
rect 935 2765 950 2785
rect 0 2750 950 2765
rect 0 2685 50 2700
rect 0 2665 15 2685
rect 35 2665 50 2685
rect 0 2635 50 2665
rect 0 2615 15 2635
rect 35 2615 50 2635
rect 0 2585 50 2615
rect 0 2565 15 2585
rect 35 2565 50 2585
rect 0 2535 50 2565
rect 0 2515 15 2535
rect 35 2515 50 2535
rect 0 2485 50 2515
rect 0 2465 15 2485
rect 35 2465 50 2485
rect 0 2435 50 2465
rect 0 2415 15 2435
rect 35 2415 50 2435
rect 0 2385 50 2415
rect 0 2365 15 2385
rect 35 2365 50 2385
rect 0 2335 50 2365
rect 0 2315 15 2335
rect 35 2315 50 2335
rect 0 2285 50 2315
rect 0 2265 15 2285
rect 35 2265 50 2285
rect 0 2235 50 2265
rect 0 2215 15 2235
rect 35 2215 50 2235
rect 0 2185 50 2215
rect 0 2165 15 2185
rect 35 2165 50 2185
rect 0 2135 50 2165
rect 0 2115 15 2135
rect 35 2115 50 2135
rect 0 2085 50 2115
rect 0 2065 15 2085
rect 35 2065 50 2085
rect 0 2035 50 2065
rect 0 2015 15 2035
rect 35 2015 50 2035
rect 0 2000 50 2015
rect 900 2685 950 2700
rect 900 2665 915 2685
rect 935 2665 950 2685
rect 900 2635 950 2665
rect 900 2615 915 2635
rect 935 2615 950 2635
rect 900 2585 950 2615
rect 900 2565 915 2585
rect 935 2565 950 2585
rect 900 2535 950 2565
rect 900 2515 915 2535
rect 935 2515 950 2535
rect 900 2485 950 2515
rect 900 2465 915 2485
rect 935 2465 950 2485
rect 900 2435 950 2465
rect 900 2415 915 2435
rect 935 2415 950 2435
rect 900 2385 950 2415
rect 900 2365 915 2385
rect 935 2365 950 2385
rect 900 2335 950 2365
rect 900 2315 915 2335
rect 935 2315 950 2335
rect 900 2285 950 2315
rect 900 2265 915 2285
rect 935 2265 950 2285
rect 900 2235 950 2265
rect 900 2215 915 2235
rect 935 2215 950 2235
rect 900 2185 950 2215
rect 900 2165 915 2185
rect 935 2165 950 2185
rect 900 2135 950 2165
rect 900 2115 915 2135
rect 935 2115 950 2135
rect 900 2085 950 2115
rect 900 2065 915 2085
rect 935 2065 950 2085
rect 900 2035 950 2065
rect 900 2015 915 2035
rect 935 2015 950 2035
rect 900 2000 950 2015
rect 50 1935 900 1950
rect 50 1915 65 1935
rect 85 1915 115 1935
rect 135 1915 165 1935
rect 185 1915 215 1935
rect 235 1915 265 1935
rect 285 1915 315 1935
rect 335 1915 365 1935
rect 385 1915 415 1935
rect 435 1915 465 1935
rect 485 1915 515 1935
rect 535 1915 565 1935
rect 585 1915 615 1935
rect 635 1915 665 1935
rect 685 1915 715 1935
rect 735 1915 765 1935
rect 785 1915 815 1935
rect 835 1915 865 1935
rect 885 1915 900 1935
rect 50 1900 900 1915
rect 0 1835 50 1850
rect 0 1815 15 1835
rect 35 1815 50 1835
rect 0 1785 50 1815
rect 0 1765 15 1785
rect 35 1765 50 1785
rect 0 1735 50 1765
rect 0 1715 15 1735
rect 35 1715 50 1735
rect 0 1685 50 1715
rect 0 1665 15 1685
rect 35 1665 50 1685
rect 0 1635 50 1665
rect 0 1615 15 1635
rect 35 1615 50 1635
rect 0 1585 50 1615
rect 0 1565 15 1585
rect 35 1565 50 1585
rect 0 1535 50 1565
rect 0 1515 15 1535
rect 35 1515 50 1535
rect 0 1485 50 1515
rect 0 1465 15 1485
rect 35 1465 50 1485
rect 0 1435 50 1465
rect 0 1415 15 1435
rect 35 1415 50 1435
rect 0 1385 50 1415
rect 0 1365 15 1385
rect 35 1365 50 1385
rect 0 1335 50 1365
rect 0 1315 15 1335
rect 35 1315 50 1335
rect 0 1285 50 1315
rect 0 1265 15 1285
rect 35 1265 50 1285
rect 0 1235 50 1265
rect 0 1215 15 1235
rect 35 1215 50 1235
rect 0 1185 50 1215
rect 0 1165 15 1185
rect 35 1165 50 1185
rect 0 1150 50 1165
rect 900 1835 950 1850
rect 900 1815 915 1835
rect 935 1815 950 1835
rect 900 1785 950 1815
rect 900 1765 915 1785
rect 935 1765 950 1785
rect 900 1735 950 1765
rect 900 1715 915 1735
rect 935 1715 950 1735
rect 900 1685 950 1715
rect 900 1665 915 1685
rect 935 1665 950 1685
rect 900 1635 950 1665
rect 900 1615 915 1635
rect 935 1615 950 1635
rect 900 1585 950 1615
rect 900 1565 915 1585
rect 935 1565 950 1585
rect 900 1535 950 1565
rect 900 1515 915 1535
rect 935 1515 950 1535
rect 900 1485 950 1515
rect 900 1465 915 1485
rect 935 1465 950 1485
rect 900 1435 950 1465
rect 900 1415 915 1435
rect 935 1415 950 1435
rect 900 1385 950 1415
rect 900 1365 915 1385
rect 935 1365 950 1385
rect 900 1335 950 1365
rect 900 1315 915 1335
rect 935 1315 950 1335
rect 900 1285 950 1315
rect 900 1265 915 1285
rect 935 1265 950 1285
rect 900 1235 950 1265
rect 900 1215 915 1235
rect 935 1215 950 1235
rect 900 1185 950 1215
rect 900 1165 915 1185
rect 935 1165 950 1185
rect 900 1150 950 1165
rect 0 1085 950 1100
rect 0 1065 15 1085
rect 35 1065 65 1085
rect 85 1065 115 1085
rect 135 1065 165 1085
rect 185 1065 215 1085
rect 235 1065 265 1085
rect 285 1065 315 1085
rect 335 1065 365 1085
rect 385 1065 415 1085
rect 435 1065 465 1085
rect 485 1065 515 1085
rect 535 1065 565 1085
rect 585 1065 615 1085
rect 635 1065 665 1085
rect 685 1065 715 1085
rect 735 1065 765 1085
rect 785 1065 815 1085
rect 835 1065 865 1085
rect 885 1065 915 1085
rect 935 1065 950 1085
rect 0 1050 950 1065
rect 0 935 950 950
rect 0 915 15 935
rect 35 915 65 935
rect 85 915 115 935
rect 135 915 165 935
rect 185 915 215 935
rect 235 915 265 935
rect 285 915 315 935
rect 335 915 365 935
rect 385 915 415 935
rect 435 915 465 935
rect 485 915 515 935
rect 535 915 565 935
rect 585 915 615 935
rect 635 915 665 935
rect 685 915 715 935
rect 735 915 765 935
rect 785 915 815 935
rect 835 915 865 935
rect 885 915 915 935
rect 935 915 950 935
rect 0 900 950 915
rect 50 835 900 850
rect 50 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 215 835
rect 235 815 265 835
rect 285 815 315 835
rect 335 815 365 835
rect 385 815 415 835
rect 435 815 465 835
rect 485 815 515 835
rect 535 815 565 835
rect 585 815 615 835
rect 635 815 665 835
rect 685 815 715 835
rect 735 815 765 835
rect 785 815 815 835
rect 835 815 865 835
rect 885 815 900 835
rect 50 800 900 815
rect 0 735 50 750
rect 0 715 15 735
rect 35 715 50 735
rect 0 685 50 715
rect 0 665 15 685
rect 35 665 50 685
rect 0 635 50 665
rect 0 615 15 635
rect 35 615 50 635
rect 0 585 50 615
rect 0 565 15 585
rect 35 565 50 585
rect 0 535 50 565
rect 0 515 15 535
rect 35 515 50 535
rect 0 485 50 515
rect 0 465 15 485
rect 35 465 50 485
rect 0 435 50 465
rect 0 415 15 435
rect 35 415 50 435
rect 0 385 50 415
rect 0 365 15 385
rect 35 365 50 385
rect 0 335 50 365
rect 0 315 15 335
rect 35 315 50 335
rect 0 285 50 315
rect 0 265 15 285
rect 35 265 50 285
rect 0 250 50 265
rect 450 735 500 750
rect 450 715 465 735
rect 485 715 500 735
rect 450 685 500 715
rect 450 665 465 685
rect 485 665 500 685
rect 450 635 500 665
rect 450 615 465 635
rect 485 615 500 635
rect 450 585 500 615
rect 450 565 465 585
rect 485 565 500 585
rect 450 535 500 565
rect 450 515 465 535
rect 485 515 500 535
rect 450 485 500 515
rect 450 465 465 485
rect 485 465 500 485
rect 450 435 500 465
rect 450 415 465 435
rect 485 415 500 435
rect 450 385 500 415
rect 450 365 465 385
rect 485 365 500 385
rect 450 335 500 365
rect 450 315 465 335
rect 485 315 500 335
rect 450 285 500 315
rect 450 265 465 285
rect 485 265 500 285
rect 450 250 500 265
rect 900 735 950 750
rect 900 715 915 735
rect 935 715 950 735
rect 900 685 950 715
rect 900 665 915 685
rect 935 665 950 685
rect 900 635 950 665
rect 900 615 915 635
rect 935 615 950 635
rect 900 585 950 615
rect 900 565 915 585
rect 935 565 950 585
rect 900 535 950 565
rect 900 515 915 535
rect 935 515 950 535
rect 900 485 950 515
rect 900 465 915 485
rect 935 465 950 485
rect 900 435 950 465
rect 900 415 915 435
rect 935 415 950 435
rect 900 385 950 415
rect 900 365 915 385
rect 935 365 950 385
rect 900 335 950 365
rect 900 315 915 335
rect 935 315 950 335
rect 900 285 950 315
rect 900 265 915 285
rect 935 265 950 285
rect 900 250 950 265
rect 0 185 950 200
rect 0 165 15 185
rect 35 165 65 185
rect 85 165 115 185
rect 135 165 165 185
rect 185 165 215 185
rect 235 165 265 185
rect 285 165 315 185
rect 335 165 365 185
rect 385 165 415 185
rect 435 165 465 185
rect 485 165 515 185
rect 535 165 565 185
rect 585 165 615 185
rect 635 165 665 185
rect 685 165 715 185
rect 735 165 765 185
rect 785 165 815 185
rect 835 165 865 185
rect 885 165 915 185
rect 935 165 950 185
rect 0 150 950 165
rect 0 35 950 50
rect 0 15 15 35
rect 35 15 65 35
rect 85 15 115 35
rect 135 15 165 35
rect 185 15 215 35
rect 235 15 265 35
rect 285 15 315 35
rect 335 15 365 35
rect 385 15 415 35
rect 435 15 465 35
rect 485 15 515 35
rect 535 15 565 35
rect 585 15 615 35
rect 635 15 665 35
rect 685 15 715 35
rect 735 15 765 35
rect 785 15 815 35
rect 835 15 865 35
rect 885 15 915 35
rect 935 15 950 35
rect 0 0 950 15
<< viali >>
rect 15 3565 35 3585
rect 15 3515 35 3535
rect 15 3465 35 3485
rect 15 3415 35 3435
rect 15 3365 35 3385
rect 15 3315 35 3335
rect 15 3265 35 3285
rect 15 3215 35 3235
rect 15 3165 35 3185
rect 15 3115 35 3135
rect 465 3565 485 3585
rect 465 3515 485 3535
rect 465 3465 485 3485
rect 465 3415 485 3435
rect 465 3365 485 3385
rect 465 3315 485 3335
rect 465 3265 485 3285
rect 465 3215 485 3235
rect 465 3165 485 3185
rect 465 3115 485 3135
rect 915 3565 935 3585
rect 915 3515 935 3535
rect 915 3465 935 3485
rect 915 3415 935 3435
rect 915 3365 935 3385
rect 915 3315 935 3335
rect 915 3265 935 3285
rect 915 3215 935 3235
rect 465 3015 485 3035
rect 15 2665 35 2685
rect 15 2615 35 2635
rect 15 2565 35 2585
rect 15 2515 35 2535
rect 15 2465 35 2485
rect 15 2415 35 2435
rect 15 2365 35 2385
rect 15 2315 35 2335
rect 15 2265 35 2285
rect 15 2215 35 2235
rect 15 2165 35 2185
rect 15 2115 35 2135
rect 15 2065 35 2085
rect 15 2015 35 2035
rect 915 2665 935 2685
rect 915 2615 935 2635
rect 915 2565 935 2585
rect 915 2515 935 2535
rect 915 2465 935 2485
rect 915 2415 935 2435
rect 915 2365 935 2385
rect 915 2315 935 2335
rect 915 2265 935 2285
rect 915 2215 935 2235
rect 915 2165 935 2185
rect 915 2115 935 2135
rect 915 2065 935 2085
rect 915 2015 935 2035
rect 465 1915 485 1935
rect 15 1815 35 1835
rect 15 1765 35 1785
rect 15 1715 35 1735
rect 15 1665 35 1685
rect 15 1615 35 1635
rect 15 1565 35 1585
rect 15 1515 35 1535
rect 15 1465 35 1485
rect 15 1415 35 1435
rect 15 1365 35 1385
rect 15 1315 35 1335
rect 15 1265 35 1285
rect 15 1215 35 1235
rect 15 1165 35 1185
rect 915 1815 935 1835
rect 915 1765 935 1785
rect 915 1715 935 1735
rect 915 1665 935 1685
rect 915 1615 935 1635
rect 915 1565 935 1585
rect 915 1515 935 1535
rect 915 1465 935 1485
rect 915 1415 935 1435
rect 915 1365 935 1385
rect 915 1315 935 1335
rect 915 1265 935 1285
rect 915 1215 935 1235
rect 915 1165 935 1185
rect 465 815 485 835
rect 15 715 35 735
rect 15 665 35 685
rect 15 615 35 635
rect 15 565 35 585
rect 15 515 35 535
rect 15 465 35 485
rect 15 415 35 435
rect 15 365 35 385
rect 15 315 35 335
rect 15 265 35 285
rect 465 715 485 735
rect 465 665 485 685
rect 465 615 485 635
rect 465 565 485 585
rect 465 515 485 535
rect 465 465 485 485
rect 465 415 485 435
rect 465 365 485 385
rect 465 315 485 335
rect 465 265 485 285
rect 915 615 935 635
rect 915 565 935 585
rect 915 515 935 535
rect 915 465 935 485
rect 915 415 935 435
rect 915 365 935 385
rect 915 315 935 335
rect 915 265 935 285
<< metal1 >>
rect 0 3740 50 3750
rect 0 3710 10 3740
rect 40 3710 50 3740
rect 0 3640 50 3710
rect 0 3610 10 3640
rect 40 3610 50 3640
rect 0 3585 50 3610
rect 900 3740 950 3750
rect 900 3710 910 3740
rect 940 3710 950 3740
rect 900 3640 950 3710
rect 900 3610 910 3640
rect 940 3610 950 3640
rect 0 3565 15 3585
rect 35 3565 50 3585
rect 0 3540 50 3565
rect 0 3510 10 3540
rect 40 3510 50 3540
rect 0 3485 50 3510
rect 0 3465 15 3485
rect 35 3465 50 3485
rect 0 3440 50 3465
rect 0 3410 10 3440
rect 40 3410 50 3440
rect 0 3385 50 3410
rect 0 3365 15 3385
rect 35 3365 50 3385
rect 0 3340 50 3365
rect 0 3310 10 3340
rect 40 3310 50 3340
rect 0 3285 50 3310
rect 0 3265 15 3285
rect 35 3265 50 3285
rect 0 3240 50 3265
rect 0 3210 10 3240
rect 40 3210 50 3240
rect 0 3185 50 3210
rect 0 3165 15 3185
rect 35 3165 50 3185
rect 0 3140 50 3165
rect 0 3110 10 3140
rect 40 3110 50 3140
rect 0 3100 50 3110
rect 450 3585 500 3600
rect 450 3565 465 3585
rect 485 3565 500 3585
rect 450 3535 500 3565
rect 450 3515 465 3535
rect 485 3515 500 3535
rect 450 3485 500 3515
rect 450 3465 465 3485
rect 485 3465 500 3485
rect 450 3435 500 3465
rect 450 3415 465 3435
rect 485 3415 500 3435
rect 450 3385 500 3415
rect 450 3365 465 3385
rect 485 3365 500 3385
rect 450 3335 500 3365
rect 450 3315 465 3335
rect 485 3315 500 3335
rect 450 3285 500 3315
rect 450 3265 465 3285
rect 485 3265 500 3285
rect 450 3235 500 3265
rect 450 3215 465 3235
rect 485 3215 500 3235
rect 450 3185 500 3215
rect 900 3585 950 3610
rect 900 3565 915 3585
rect 935 3565 950 3585
rect 900 3540 950 3565
rect 900 3510 910 3540
rect 940 3510 950 3540
rect 900 3485 950 3510
rect 900 3465 915 3485
rect 935 3465 950 3485
rect 900 3440 950 3465
rect 900 3410 910 3440
rect 940 3410 950 3440
rect 900 3385 950 3410
rect 900 3365 915 3385
rect 935 3365 950 3385
rect 900 3340 950 3365
rect 900 3310 910 3340
rect 940 3310 950 3340
rect 900 3285 950 3310
rect 900 3265 915 3285
rect 935 3265 950 3285
rect 900 3240 950 3265
rect 900 3210 910 3240
rect 940 3210 950 3240
rect 900 3200 950 3210
rect 450 3165 465 3185
rect 485 3165 500 3185
rect 450 3150 500 3165
rect 450 3135 950 3150
rect 450 3115 465 3135
rect 485 3115 950 3135
rect 450 3100 950 3115
rect 450 3040 500 3050
rect 450 3010 460 3040
rect 490 3010 500 3040
rect 450 3000 500 3010
rect 0 2840 50 2850
rect 0 2810 10 2840
rect 40 2810 50 2840
rect 0 2685 50 2810
rect 0 2665 15 2685
rect 35 2665 50 2685
rect 0 2635 50 2665
rect 0 2615 15 2635
rect 35 2615 50 2635
rect 0 2585 50 2615
rect 0 2565 15 2585
rect 35 2565 50 2585
rect 0 2535 50 2565
rect 0 2515 15 2535
rect 35 2515 50 2535
rect 0 2485 50 2515
rect 0 2465 15 2485
rect 35 2465 50 2485
rect 0 2440 50 2465
rect 0 2410 10 2440
rect 40 2410 50 2440
rect 0 2385 50 2410
rect 0 2365 15 2385
rect 35 2365 50 2385
rect 0 2335 50 2365
rect 0 2315 15 2335
rect 35 2315 50 2335
rect 0 2285 50 2315
rect 0 2265 15 2285
rect 35 2265 50 2285
rect 0 2240 50 2265
rect 0 2210 10 2240
rect 40 2210 50 2240
rect 0 2185 50 2210
rect 0 2165 15 2185
rect 35 2165 50 2185
rect 0 2135 50 2165
rect 0 2115 15 2135
rect 35 2115 50 2135
rect 0 2085 50 2115
rect 0 2065 15 2085
rect 35 2065 50 2085
rect 0 2040 50 2065
rect 0 2010 10 2040
rect 40 2010 50 2040
rect 0 1840 50 2010
rect 900 2685 950 3100
rect 900 2665 915 2685
rect 935 2665 950 2685
rect 900 2635 950 2665
rect 900 2615 915 2635
rect 935 2615 950 2635
rect 900 2585 950 2615
rect 900 2565 915 2585
rect 935 2565 950 2585
rect 900 2535 950 2565
rect 900 2515 915 2535
rect 935 2515 950 2535
rect 900 2485 950 2515
rect 900 2465 915 2485
rect 935 2465 950 2485
rect 900 2435 950 2465
rect 900 2415 915 2435
rect 935 2415 950 2435
rect 900 2385 950 2415
rect 900 2365 915 2385
rect 935 2365 950 2385
rect 900 2335 950 2365
rect 900 2315 915 2335
rect 935 2315 950 2335
rect 900 2285 950 2315
rect 900 2265 915 2285
rect 935 2265 950 2285
rect 900 2235 950 2265
rect 900 2215 915 2235
rect 935 2215 950 2235
rect 900 2185 950 2215
rect 900 2165 915 2185
rect 935 2165 950 2185
rect 900 2135 950 2165
rect 900 2115 915 2135
rect 935 2115 950 2135
rect 900 2085 950 2115
rect 900 2065 915 2085
rect 935 2065 950 2085
rect 900 2035 950 2065
rect 900 2015 915 2035
rect 935 2015 950 2035
rect 450 1940 500 1950
rect 450 1910 460 1940
rect 490 1910 500 1940
rect 450 1900 500 1910
rect 0 1810 10 1840
rect 40 1810 50 1840
rect 0 1785 50 1810
rect 0 1765 15 1785
rect 35 1765 50 1785
rect 0 1735 50 1765
rect 0 1715 15 1735
rect 35 1715 50 1735
rect 0 1685 50 1715
rect 0 1665 15 1685
rect 35 1665 50 1685
rect 0 1640 50 1665
rect 0 1610 10 1640
rect 40 1610 50 1640
rect 0 1585 50 1610
rect 0 1565 15 1585
rect 35 1565 50 1585
rect 0 1535 50 1565
rect 0 1515 15 1535
rect 35 1515 50 1535
rect 0 1485 50 1515
rect 0 1465 15 1485
rect 35 1465 50 1485
rect 0 1440 50 1465
rect 0 1410 10 1440
rect 40 1410 50 1440
rect 0 1385 50 1410
rect 0 1365 15 1385
rect 35 1365 50 1385
rect 0 1335 50 1365
rect 0 1315 15 1335
rect 35 1315 50 1335
rect 0 1285 50 1315
rect 0 1265 15 1285
rect 35 1265 50 1285
rect 0 1235 50 1265
rect 0 1215 15 1235
rect 35 1215 50 1235
rect 0 1185 50 1215
rect 0 1165 15 1185
rect 35 1165 50 1185
rect 0 1040 50 1165
rect 0 1010 10 1040
rect 40 1010 50 1040
rect 0 1000 50 1010
rect 900 1835 950 2015
rect 900 1815 915 1835
rect 935 1815 950 1835
rect 900 1785 950 1815
rect 900 1765 915 1785
rect 935 1765 950 1785
rect 900 1735 950 1765
rect 900 1715 915 1735
rect 935 1715 950 1735
rect 900 1685 950 1715
rect 900 1665 915 1685
rect 935 1665 950 1685
rect 900 1635 950 1665
rect 900 1615 915 1635
rect 935 1615 950 1635
rect 900 1585 950 1615
rect 900 1565 915 1585
rect 935 1565 950 1585
rect 900 1535 950 1565
rect 900 1515 915 1535
rect 935 1515 950 1535
rect 900 1485 950 1515
rect 900 1465 915 1485
rect 935 1465 950 1485
rect 900 1435 950 1465
rect 900 1415 915 1435
rect 935 1415 950 1435
rect 900 1385 950 1415
rect 900 1365 915 1385
rect 935 1365 950 1385
rect 900 1335 950 1365
rect 900 1315 915 1335
rect 935 1315 950 1335
rect 900 1285 950 1315
rect 900 1265 915 1285
rect 935 1265 950 1285
rect 900 1235 950 1265
rect 900 1215 915 1235
rect 935 1215 950 1235
rect 900 1185 950 1215
rect 900 1165 915 1185
rect 935 1165 950 1185
rect 450 840 500 850
rect 450 810 460 840
rect 490 810 500 840
rect 450 800 500 810
rect 900 750 950 1165
rect 0 740 50 750
rect 0 710 10 740
rect 40 710 50 740
rect 0 685 50 710
rect 0 665 15 685
rect 35 665 50 685
rect 0 640 50 665
rect 0 610 10 640
rect 40 610 50 640
rect 0 585 50 610
rect 0 565 15 585
rect 35 565 50 585
rect 0 540 50 565
rect 0 510 10 540
rect 40 510 50 540
rect 0 485 50 510
rect 0 465 15 485
rect 35 465 50 485
rect 0 440 50 465
rect 0 410 10 440
rect 40 410 50 440
rect 0 385 50 410
rect 0 365 15 385
rect 35 365 50 385
rect 0 340 50 365
rect 0 310 10 340
rect 40 310 50 340
rect 0 285 50 310
rect 0 265 15 285
rect 35 265 50 285
rect 0 240 50 265
rect 450 735 950 750
rect 450 715 465 735
rect 485 715 950 735
rect 450 700 950 715
rect 450 685 500 700
rect 450 665 465 685
rect 485 665 500 685
rect 450 635 500 665
rect 450 615 465 635
rect 485 615 500 635
rect 450 585 500 615
rect 450 565 465 585
rect 485 565 500 585
rect 450 535 500 565
rect 450 515 465 535
rect 485 515 500 535
rect 450 485 500 515
rect 450 465 465 485
rect 485 465 500 485
rect 450 435 500 465
rect 450 415 465 435
rect 485 415 500 435
rect 450 385 500 415
rect 450 365 465 385
rect 485 365 500 385
rect 450 335 500 365
rect 450 315 465 335
rect 485 315 500 335
rect 450 285 500 315
rect 450 265 465 285
rect 485 265 500 285
rect 450 250 500 265
rect 900 640 950 650
rect 900 610 910 640
rect 940 610 950 640
rect 900 585 950 610
rect 900 565 915 585
rect 935 565 950 585
rect 900 540 950 565
rect 900 510 910 540
rect 940 510 950 540
rect 900 485 950 510
rect 900 465 915 485
rect 935 465 950 485
rect 900 440 950 465
rect 900 410 910 440
rect 940 410 950 440
rect 900 385 950 410
rect 900 365 915 385
rect 935 365 950 385
rect 900 340 950 365
rect 900 310 910 340
rect 940 310 950 340
rect 900 285 950 310
rect 900 265 915 285
rect 935 265 950 285
rect 0 210 10 240
rect 40 210 50 240
rect 0 140 50 210
rect 0 110 10 140
rect 40 110 50 140
rect 0 100 50 110
rect 900 240 950 265
rect 900 210 910 240
rect 940 210 950 240
rect 900 140 950 210
rect 900 110 910 140
rect 940 110 950 140
rect 900 100 950 110
<< via1 >>
rect 10 3710 40 3740
rect 10 3610 40 3640
rect 910 3710 940 3740
rect 910 3610 940 3640
rect 10 3535 40 3540
rect 10 3515 15 3535
rect 15 3515 35 3535
rect 35 3515 40 3535
rect 10 3510 40 3515
rect 10 3435 40 3440
rect 10 3415 15 3435
rect 15 3415 35 3435
rect 35 3415 40 3435
rect 10 3410 40 3415
rect 10 3335 40 3340
rect 10 3315 15 3335
rect 15 3315 35 3335
rect 35 3315 40 3335
rect 10 3310 40 3315
rect 10 3235 40 3240
rect 10 3215 15 3235
rect 15 3215 35 3235
rect 35 3215 40 3235
rect 10 3210 40 3215
rect 10 3135 40 3140
rect 10 3115 15 3135
rect 15 3115 35 3135
rect 35 3115 40 3135
rect 10 3110 40 3115
rect 910 3535 940 3540
rect 910 3515 915 3535
rect 915 3515 935 3535
rect 935 3515 940 3535
rect 910 3510 940 3515
rect 910 3435 940 3440
rect 910 3415 915 3435
rect 915 3415 935 3435
rect 935 3415 940 3435
rect 910 3410 940 3415
rect 910 3335 940 3340
rect 910 3315 915 3335
rect 915 3315 935 3335
rect 935 3315 940 3335
rect 910 3310 940 3315
rect 910 3235 940 3240
rect 910 3215 915 3235
rect 915 3215 935 3235
rect 935 3215 940 3235
rect 910 3210 940 3215
rect 460 3035 490 3040
rect 460 3015 465 3035
rect 465 3015 485 3035
rect 485 3015 490 3035
rect 460 3010 490 3015
rect 10 2810 40 2840
rect 10 2435 40 2440
rect 10 2415 15 2435
rect 15 2415 35 2435
rect 35 2415 40 2435
rect 10 2410 40 2415
rect 10 2235 40 2240
rect 10 2215 15 2235
rect 15 2215 35 2235
rect 35 2215 40 2235
rect 10 2210 40 2215
rect 10 2035 40 2040
rect 10 2015 15 2035
rect 15 2015 35 2035
rect 35 2015 40 2035
rect 10 2010 40 2015
rect 460 1935 490 1940
rect 460 1915 465 1935
rect 465 1915 485 1935
rect 485 1915 490 1935
rect 460 1910 490 1915
rect 10 1835 40 1840
rect 10 1815 15 1835
rect 15 1815 35 1835
rect 35 1815 40 1835
rect 10 1810 40 1815
rect 10 1635 40 1640
rect 10 1615 15 1635
rect 15 1615 35 1635
rect 35 1615 40 1635
rect 10 1610 40 1615
rect 10 1435 40 1440
rect 10 1415 15 1435
rect 15 1415 35 1435
rect 35 1415 40 1435
rect 10 1410 40 1415
rect 10 1010 40 1040
rect 460 835 490 840
rect 460 815 465 835
rect 465 815 485 835
rect 485 815 490 835
rect 460 810 490 815
rect 10 735 40 740
rect 10 715 15 735
rect 15 715 35 735
rect 35 715 40 735
rect 10 710 40 715
rect 10 635 40 640
rect 10 615 15 635
rect 15 615 35 635
rect 35 615 40 635
rect 10 610 40 615
rect 10 535 40 540
rect 10 515 15 535
rect 15 515 35 535
rect 35 515 40 535
rect 10 510 40 515
rect 10 435 40 440
rect 10 415 15 435
rect 15 415 35 435
rect 35 415 40 435
rect 10 410 40 415
rect 10 335 40 340
rect 10 315 15 335
rect 15 315 35 335
rect 35 315 40 335
rect 10 310 40 315
rect 910 635 940 640
rect 910 615 915 635
rect 915 615 935 635
rect 935 615 940 635
rect 910 610 940 615
rect 910 535 940 540
rect 910 515 915 535
rect 915 515 935 535
rect 935 515 940 535
rect 910 510 940 515
rect 910 435 940 440
rect 910 415 915 435
rect 915 415 935 435
rect 935 415 940 435
rect 910 410 940 415
rect 910 335 940 340
rect 910 315 915 335
rect 915 315 935 335
rect 935 315 940 335
rect 910 310 940 315
rect 10 210 40 240
rect 10 110 40 140
rect 910 210 940 240
rect 910 110 940 140
<< metal2 >>
rect 0 3740 950 3750
rect 0 3710 10 3740
rect 40 3710 910 3740
rect 940 3710 950 3740
rect 0 3700 950 3710
rect 0 3640 950 3650
rect 0 3610 10 3640
rect 40 3610 910 3640
rect 940 3610 950 3640
rect 0 3600 950 3610
rect 0 3540 950 3550
rect 0 3510 10 3540
rect 40 3510 910 3540
rect 940 3510 950 3540
rect 0 3500 950 3510
rect 0 3440 950 3450
rect 0 3410 10 3440
rect 40 3410 910 3440
rect 940 3410 950 3440
rect 0 3400 950 3410
rect 0 3340 950 3350
rect 0 3310 10 3340
rect 40 3310 910 3340
rect 940 3310 950 3340
rect 0 3300 950 3310
rect 0 3240 950 3250
rect 0 3210 10 3240
rect 40 3210 910 3240
rect 940 3210 950 3240
rect 0 3200 950 3210
rect 0 3140 950 3150
rect 0 3110 10 3140
rect 40 3110 910 3140
rect 940 3110 950 3140
rect 0 3100 950 3110
rect 450 3040 500 3050
rect 450 3010 460 3040
rect 490 3010 500 3040
rect 450 3000 500 3010
rect 0 2840 950 2850
rect 0 2810 10 2840
rect 40 2810 910 2840
rect 940 2810 950 2840
rect 0 2800 950 2810
rect 0 2440 950 2450
rect 0 2410 10 2440
rect 40 2410 950 2440
rect 0 2400 950 2410
rect 0 2240 950 2250
rect 0 2210 10 2240
rect 40 2210 950 2240
rect 0 2200 950 2210
rect 0 2040 950 2050
rect 0 2010 10 2040
rect 40 2010 950 2040
rect 0 2000 950 2010
rect 450 1940 500 1950
rect 450 1910 460 1940
rect 490 1910 500 1940
rect 450 1900 500 1910
rect 0 1840 950 1850
rect 0 1810 10 1840
rect 40 1810 950 1840
rect 0 1800 950 1810
rect 0 1640 950 1650
rect 0 1610 10 1640
rect 40 1610 950 1640
rect 0 1600 950 1610
rect 0 1440 950 1450
rect 0 1410 10 1440
rect 40 1410 950 1440
rect 0 1400 950 1410
rect 0 1040 950 1050
rect 0 1010 10 1040
rect 40 1010 910 1040
rect 940 1010 950 1040
rect 0 1000 950 1010
rect 450 840 500 850
rect 450 810 460 840
rect 490 810 500 840
rect 450 800 500 810
rect 0 740 950 750
rect 0 710 10 740
rect 40 710 910 740
rect 940 710 950 740
rect 0 700 950 710
rect 0 640 950 650
rect 0 610 10 640
rect 40 610 910 640
rect 940 610 950 640
rect 0 600 950 610
rect 450 550 500 600
rect 0 540 950 550
rect 0 510 10 540
rect 40 510 910 540
rect 940 510 950 540
rect 0 500 950 510
rect 450 450 500 500
rect 0 440 950 450
rect 0 410 10 440
rect 40 410 910 440
rect 940 410 950 440
rect 0 400 950 410
rect 450 350 500 400
rect 0 340 950 350
rect 0 310 10 340
rect 40 310 910 340
rect 940 310 950 340
rect 0 300 950 310
rect 450 250 500 300
rect 0 240 950 250
rect 0 210 10 240
rect 40 210 910 240
rect 940 210 950 240
rect 0 200 950 210
rect 0 140 950 150
rect 0 110 10 140
rect 40 110 910 140
rect 940 110 950 140
rect 0 100 950 110
<< via2 >>
rect 10 3710 40 3740
rect 910 3710 940 3740
rect 10 3610 40 3640
rect 910 3610 940 3640
rect 10 3510 40 3540
rect 910 3510 940 3540
rect 10 3410 40 3440
rect 910 3410 940 3440
rect 10 3310 40 3340
rect 910 3310 940 3340
rect 10 3210 40 3240
rect 910 3210 940 3240
rect 10 3110 40 3140
rect 910 3110 940 3140
rect 460 3010 490 3040
rect 10 2810 40 2840
rect 910 2810 940 2840
rect 10 2410 40 2440
rect 10 2210 40 2240
rect 10 2010 40 2040
rect 460 1910 490 1940
rect 10 1810 40 1840
rect 10 1610 40 1640
rect 10 1410 40 1440
rect 10 1010 40 1040
rect 910 1010 940 1040
rect 460 810 490 840
rect 10 710 40 740
rect 910 710 940 740
rect 10 610 40 640
rect 910 610 940 640
rect 10 510 40 540
rect 910 510 940 540
rect 10 410 40 440
rect 910 410 940 440
rect 10 310 40 340
rect 910 310 940 340
rect 10 210 40 240
rect 910 210 940 240
rect 10 110 40 140
rect 910 110 940 140
<< metal3 >>
rect 0 3740 950 3750
rect 0 3710 10 3740
rect 40 3710 910 3740
rect 940 3710 950 3740
rect 0 3700 950 3710
rect 0 3640 950 3650
rect 0 3610 10 3640
rect 40 3610 910 3640
rect 940 3610 950 3640
rect 0 3600 950 3610
rect 0 3540 950 3550
rect 0 3510 10 3540
rect 40 3510 910 3540
rect 940 3510 950 3540
rect 0 3500 950 3510
rect 0 3440 950 3450
rect 0 3410 10 3440
rect 40 3410 910 3440
rect 940 3410 950 3440
rect 0 3400 950 3410
rect 0 3340 950 3350
rect 0 3310 10 3340
rect 40 3310 910 3340
rect 940 3310 950 3340
rect 0 3300 950 3310
rect 0 3240 950 3250
rect 0 3210 10 3240
rect 40 3210 910 3240
rect 940 3210 950 3240
rect 0 3200 950 3210
rect 0 3140 950 3150
rect 0 3110 10 3140
rect 40 3110 910 3140
rect 940 3110 950 3140
rect 0 3100 950 3110
rect 450 3045 500 3050
rect 450 3005 455 3045
rect 495 3005 500 3045
rect 450 3000 500 3005
rect 0 2840 950 2850
rect 0 2810 10 2840
rect 40 2810 910 2840
rect 940 2810 950 2840
rect 0 2800 950 2810
rect 0 2440 950 2450
rect 0 2410 10 2440
rect 40 2410 950 2440
rect 0 2400 950 2410
rect 0 2240 950 2250
rect 0 2210 10 2240
rect 40 2210 950 2240
rect 0 2200 950 2210
rect 0 2040 950 2050
rect 0 2010 10 2040
rect 40 2010 950 2040
rect 0 2000 950 2010
rect 450 1945 500 1950
rect 450 1905 455 1945
rect 495 1905 500 1945
rect 450 1900 500 1905
rect 0 1840 950 1850
rect 0 1810 10 1840
rect 40 1810 950 1840
rect 0 1800 950 1810
rect 0 1640 950 1650
rect 0 1610 10 1640
rect 40 1610 950 1640
rect 0 1600 950 1610
rect 0 1440 950 1450
rect 0 1410 10 1440
rect 40 1410 950 1440
rect 0 1400 950 1410
rect 0 1040 950 1050
rect 0 1010 10 1040
rect 40 1010 910 1040
rect 940 1010 950 1040
rect 0 1000 950 1010
rect 450 845 500 850
rect 450 805 455 845
rect 495 805 500 845
rect 450 800 500 805
rect 0 740 950 750
rect 0 710 10 740
rect 40 710 910 740
rect 940 710 950 740
rect 0 700 950 710
rect 0 640 950 650
rect 0 610 10 640
rect 40 610 910 640
rect 940 610 950 640
rect 0 600 950 610
rect 450 550 500 600
rect 0 540 950 550
rect 0 510 10 540
rect 40 510 910 540
rect 940 510 950 540
rect 0 500 950 510
rect 450 450 500 500
rect 0 440 950 450
rect 0 410 10 440
rect 40 410 910 440
rect 940 410 950 440
rect 0 400 950 410
rect 450 350 500 400
rect 0 340 950 350
rect 0 310 10 340
rect 40 310 910 340
rect 940 310 950 340
rect 0 300 950 310
rect 450 250 500 300
rect 0 240 950 250
rect 0 210 10 240
rect 40 210 910 240
rect 940 210 950 240
rect 0 200 950 210
rect 0 140 950 150
rect 0 110 10 140
rect 40 110 910 140
rect 940 110 950 140
rect 0 100 950 110
<< via3 >>
rect 455 3040 495 3045
rect 455 3010 460 3040
rect 460 3010 490 3040
rect 490 3010 495 3040
rect 455 3005 495 3010
rect 455 1940 495 1945
rect 455 1910 460 1940
rect 460 1910 490 1940
rect 490 1910 495 1940
rect 455 1905 495 1910
rect 455 840 495 845
rect 455 810 460 840
rect 460 810 490 840
rect 490 810 495 840
rect 455 805 495 810
<< metal4 >>
rect 450 3045 500 3050
rect 450 3005 455 3045
rect 495 3005 500 3045
rect 450 1945 500 3005
rect 450 1905 455 1945
rect 495 1905 500 1945
rect 450 845 500 1905
rect 450 805 455 845
rect 495 805 500 845
rect 450 800 500 805
<< labels >>
rlabel metal4 450 1900 500 1950 0 in
port 1 nsew
rlabel metal1 900 1900 950 1950 0 out
port 2 nsew
rlabel locali 0 2900 950 2950 0 bp
port 3 nsew
rlabel locali 0 900 950 950 0 bp
port 3 nsew
rlabel locali 0 2750 950 2800 0 bn
port 4 nsew
rlabel locali 0 1050 950 1100 0 bn
port 4 nsew
rlabel metal3 0 3700 950 3750 0 vreg
port 5 nsew
rlabel metal3 0 100 950 150 0 vreg
port 5 nsew
rlabel metal3 0 2800 950 2850 0 vss
port 6 nsew
rlabel metal3 0 1000 950 1050 0 vss
port 6 nsew
rlabel locali 0 3800 950 3850 0 vsub
port 7 nsew
rlabel locali 0 0 950 50 0 vsub
port 7 nsew
rlabel ndiff 450 2050 500 2700 0 xt
rlabel ndiff 450 1150 500 1800 0 xb
<< end >>
