magic
tech sky130A
timestamp 1726445930
<< locali >>
rect 50 3800 3700 3850
rect 50 2900 3700 2950
rect 50 2750 3700 2800
rect 2750 2535 2800 2550
rect 2750 2515 2765 2535
rect 2785 2515 2800 2535
rect 2750 2500 2800 2515
rect 50 1050 3700 1100
rect 50 900 3700 950
rect 50 0 3700 50
<< viali >>
rect 2765 2515 2785 2535
<< metal1 >>
rect 2750 2740 2800 2750
rect 2750 2710 2760 2740
rect 2790 2710 2800 2740
rect 2750 2700 2800 2710
rect 2750 2540 2800 2550
rect 2750 2510 2760 2540
rect 2790 2510 2800 2540
rect 2750 2500 2800 2510
rect 950 1140 1000 1150
rect 950 1110 960 1140
rect 990 1110 1000 1140
rect 950 1100 1000 1110
<< via1 >>
rect 2760 2710 2790 2740
rect 2760 2510 2790 2540
rect 960 1310 990 1340
rect 960 1110 990 1140
<< metal2 >>
rect 2750 2740 2800 2750
rect 2750 2710 2760 2740
rect 2790 2710 2800 2740
rect 2750 2700 2800 2710
rect 2750 2540 2800 2550
rect 2750 2510 2760 2540
rect 2790 2510 2800 2540
rect 2750 2500 2800 2510
rect 950 1340 1000 1350
rect 950 1310 960 1340
rect 990 1310 1000 1340
rect 950 1300 1000 1310
rect 950 1140 1000 1150
rect 950 1110 960 1140
rect 990 1110 1000 1140
rect 950 1100 1000 1110
<< via2 >>
rect 2760 2710 2790 2740
rect 2760 2510 2790 2540
rect 960 1310 990 1340
rect 960 1110 990 1140
<< metal3 >>
rect 50 3700 3700 3750
rect 50 2800 3700 2850
rect 50 2740 3700 2750
rect 50 2710 2760 2740
rect 2790 2710 3700 2740
rect 50 2700 3700 2710
rect 50 2645 3700 2650
rect 50 2605 2305 2645
rect 2345 2605 3700 2645
rect 50 2600 3700 2605
rect 50 2540 3700 2550
rect 50 2510 2760 2540
rect 2790 2510 3700 2540
rect 50 2500 3700 2510
rect 50 2145 3700 2150
rect 50 2105 505 2145
rect 545 2105 3700 2145
rect 50 2100 3700 2105
rect 50 1745 3700 1750
rect 50 1705 3205 1745
rect 3245 1705 3700 1745
rect 50 1700 3700 1705
rect 50 1340 3700 1350
rect 50 1310 960 1340
rect 990 1310 3700 1340
rect 50 1300 3700 1310
rect 50 1245 3700 1250
rect 50 1205 1405 1245
rect 1445 1205 3700 1245
rect 50 1200 3700 1205
rect 50 1140 3700 1150
rect 50 1110 960 1140
rect 990 1110 3700 1140
rect 50 1100 3700 1110
rect 50 1000 3700 1050
rect 50 100 3700 150
<< via3 >>
rect 2305 2605 2345 2645
rect 505 2105 545 2145
rect 3205 1705 3245 1745
rect 1405 1205 1445 1245
<< metal4 >>
rect 2300 2645 2350 2650
rect 2300 2605 2305 2645
rect 2345 2605 2350 2645
rect 2300 2600 2350 2605
rect 500 2145 550 2150
rect 500 2105 505 2145
rect 545 2105 550 2145
rect 500 2100 550 2105
rect 3200 1745 3250 1750
rect 3200 1705 3205 1745
rect 3245 1705 3250 1745
rect 3200 1700 3250 1705
rect 1400 1245 1450 1250
rect 1400 1205 1405 1245
rect 1445 1205 1450 1245
rect 1400 1200 1450 1205
use inv1p1  a0
timestamp 1726000395
transform 1 0 50 0 1 0
box -50 0 1000 3850
use inv1p1  a1
timestamp 1726000395
transform -1 0 1900 0 1 0
box -50 0 1000 3850
use inv1p1  a2
timestamp 1726000395
transform 1 0 1850 0 1 0
box -50 0 1000 3850
use inv1p1  a3
timestamp 1726000395
transform -1 0 3700 0 1 0
box -50 0 1000 3850
<< labels >>
rlabel metal3 50 2100 3700 2150 0 ip
port 1 nsew
rlabel metal3 50 1700 3700 1750 0 im
port 2 nsew
rlabel metal3 50 2600 3700 2650 0 xm
port 3 nsew
rlabel metal3 50 1200 3700 1250 0 xp
port 4 nsew
rlabel metal3 50 2700 3700 2750 0 op
port 5 nsew
rlabel metal3 50 2500 3700 2550 0 op
port 5 nsew
rlabel metal3 50 1300 3700 1350 0 om
port 6 nsew
rlabel metal3 50 1100 3700 1150 0 om
port 6 nsew
rlabel locali 50 2900 3700 2950 0 bp
port 7 nsew
rlabel locali 50 900 3700 950 0 bp
port 7 nsew
rlabel locali 50 2750 3700 2800 0 bn
port 8 nsew
rlabel locali 50 1050 3700 1100 0 bn
port 8 nsew
rlabel metal3 50 3700 3700 3750 0 vdd
port 9 nsew
rlabel metal3 50 100 3700 150 0 vdd
port 9 nsew
rlabel metal3 50 2800 3700 2850 0 vss
port 10 nsew
rlabel metal3 50 1000 3700 1050 0 vss
port 10 nsew
rlabel locali 50 3800 3700 3850 0 vsub
port 11 nsew
rlabel locali 50 0 3700 50 0 vsub
port 11 nsew
<< end >>
