magic
tech sky130A
timestamp 1722856725
<< error_p >>
rect 250 895 300 2955
<< dnwell >>
rect 0 895 250 2955
<< nwell >>
rect -50 2850 300 3750
rect -50 100 300 1000
<< pwell >>
rect 0 1000 250 2850
<< pmoslvt >>
rect 50 3100 100 3600
rect 150 3100 200 3600
rect 50 250 100 750
rect 150 250 200 750
<< nmoslvt >>
rect 50 2000 100 2700
rect 150 2000 200 2700
rect 50 1150 100 1850
rect 150 1150 200 1850
<< ndiff >>
rect 0 2685 50 2700
rect 0 2665 15 2685
rect 35 2665 50 2685
rect 0 2635 50 2665
rect 0 2615 15 2635
rect 35 2615 50 2635
rect 0 2585 50 2615
rect 0 2565 15 2585
rect 35 2565 50 2585
rect 0 2535 50 2565
rect 0 2515 15 2535
rect 35 2515 50 2535
rect 0 2485 50 2515
rect 0 2465 15 2485
rect 35 2465 50 2485
rect 0 2435 50 2465
rect 0 2415 15 2435
rect 35 2415 50 2435
rect 0 2385 50 2415
rect 0 2365 15 2385
rect 35 2365 50 2385
rect 0 2335 50 2365
rect 0 2315 15 2335
rect 35 2315 50 2335
rect 0 2285 50 2315
rect 0 2265 15 2285
rect 35 2265 50 2285
rect 0 2235 50 2265
rect 0 2215 15 2235
rect 35 2215 50 2235
rect 0 2185 50 2215
rect 0 2165 15 2185
rect 35 2165 50 2185
rect 0 2135 50 2165
rect 0 2115 15 2135
rect 35 2115 50 2135
rect 0 2085 50 2115
rect 0 2065 15 2085
rect 35 2065 50 2085
rect 0 2035 50 2065
rect 0 2015 15 2035
rect 35 2015 50 2035
rect 0 2000 50 2015
rect 100 2685 150 2700
rect 100 2665 115 2685
rect 135 2665 150 2685
rect 100 2635 150 2665
rect 100 2615 115 2635
rect 135 2615 150 2635
rect 100 2585 150 2615
rect 100 2565 115 2585
rect 135 2565 150 2585
rect 100 2535 150 2565
rect 100 2515 115 2535
rect 135 2515 150 2535
rect 100 2485 150 2515
rect 100 2465 115 2485
rect 135 2465 150 2485
rect 100 2435 150 2465
rect 100 2415 115 2435
rect 135 2415 150 2435
rect 100 2385 150 2415
rect 100 2365 115 2385
rect 135 2365 150 2385
rect 100 2335 150 2365
rect 100 2315 115 2335
rect 135 2315 150 2335
rect 100 2285 150 2315
rect 100 2265 115 2285
rect 135 2265 150 2285
rect 100 2235 150 2265
rect 100 2215 115 2235
rect 135 2215 150 2235
rect 100 2185 150 2215
rect 100 2165 115 2185
rect 135 2165 150 2185
rect 100 2135 150 2165
rect 100 2115 115 2135
rect 135 2115 150 2135
rect 100 2085 150 2115
rect 100 2065 115 2085
rect 135 2065 150 2085
rect 100 2035 150 2065
rect 100 2015 115 2035
rect 135 2015 150 2035
rect 100 2000 150 2015
rect 200 2685 250 2700
rect 200 2665 215 2685
rect 235 2665 250 2685
rect 200 2635 250 2665
rect 200 2615 215 2635
rect 235 2615 250 2635
rect 200 2585 250 2615
rect 200 2565 215 2585
rect 235 2565 250 2585
rect 200 2535 250 2565
rect 200 2515 215 2535
rect 235 2515 250 2535
rect 200 2485 250 2515
rect 200 2465 215 2485
rect 235 2465 250 2485
rect 200 2435 250 2465
rect 200 2415 215 2435
rect 235 2415 250 2435
rect 200 2385 250 2415
rect 200 2365 215 2385
rect 235 2365 250 2385
rect 200 2335 250 2365
rect 200 2315 215 2335
rect 235 2315 250 2335
rect 200 2285 250 2315
rect 200 2265 215 2285
rect 235 2265 250 2285
rect 200 2235 250 2265
rect 200 2215 215 2235
rect 235 2215 250 2235
rect 200 2185 250 2215
rect 200 2165 215 2185
rect 235 2165 250 2185
rect 200 2135 250 2165
rect 200 2115 215 2135
rect 235 2115 250 2135
rect 200 2085 250 2115
rect 200 2065 215 2085
rect 235 2065 250 2085
rect 200 2035 250 2065
rect 200 2015 215 2035
rect 235 2015 250 2035
rect 200 2000 250 2015
rect 0 1835 50 1850
rect 0 1815 15 1835
rect 35 1815 50 1835
rect 0 1785 50 1815
rect 0 1765 15 1785
rect 35 1765 50 1785
rect 0 1735 50 1765
rect 0 1715 15 1735
rect 35 1715 50 1735
rect 0 1685 50 1715
rect 0 1665 15 1685
rect 35 1665 50 1685
rect 0 1635 50 1665
rect 0 1615 15 1635
rect 35 1615 50 1635
rect 0 1585 50 1615
rect 0 1565 15 1585
rect 35 1565 50 1585
rect 0 1535 50 1565
rect 0 1515 15 1535
rect 35 1515 50 1535
rect 0 1485 50 1515
rect 0 1465 15 1485
rect 35 1465 50 1485
rect 0 1435 50 1465
rect 0 1415 15 1435
rect 35 1415 50 1435
rect 0 1385 50 1415
rect 0 1365 15 1385
rect 35 1365 50 1385
rect 0 1335 50 1365
rect 0 1315 15 1335
rect 35 1315 50 1335
rect 0 1285 50 1315
rect 0 1265 15 1285
rect 35 1265 50 1285
rect 0 1235 50 1265
rect 0 1215 15 1235
rect 35 1215 50 1235
rect 0 1185 50 1215
rect 0 1165 15 1185
rect 35 1165 50 1185
rect 0 1150 50 1165
rect 100 1835 150 1850
rect 100 1815 115 1835
rect 135 1815 150 1835
rect 100 1785 150 1815
rect 100 1765 115 1785
rect 135 1765 150 1785
rect 100 1735 150 1765
rect 100 1715 115 1735
rect 135 1715 150 1735
rect 100 1685 150 1715
rect 100 1665 115 1685
rect 135 1665 150 1685
rect 100 1635 150 1665
rect 100 1615 115 1635
rect 135 1615 150 1635
rect 100 1585 150 1615
rect 100 1565 115 1585
rect 135 1565 150 1585
rect 100 1535 150 1565
rect 100 1515 115 1535
rect 135 1515 150 1535
rect 100 1485 150 1515
rect 100 1465 115 1485
rect 135 1465 150 1485
rect 100 1435 150 1465
rect 100 1415 115 1435
rect 135 1415 150 1435
rect 100 1385 150 1415
rect 100 1365 115 1385
rect 135 1365 150 1385
rect 100 1335 150 1365
rect 100 1315 115 1335
rect 135 1315 150 1335
rect 100 1285 150 1315
rect 100 1265 115 1285
rect 135 1265 150 1285
rect 100 1235 150 1265
rect 100 1215 115 1235
rect 135 1215 150 1235
rect 100 1185 150 1215
rect 100 1165 115 1185
rect 135 1165 150 1185
rect 100 1150 150 1165
rect 200 1835 250 1850
rect 200 1815 215 1835
rect 235 1815 250 1835
rect 200 1785 250 1815
rect 200 1765 215 1785
rect 235 1765 250 1785
rect 200 1735 250 1765
rect 200 1715 215 1735
rect 235 1715 250 1735
rect 200 1685 250 1715
rect 200 1665 215 1685
rect 235 1665 250 1685
rect 200 1635 250 1665
rect 200 1615 215 1635
rect 235 1615 250 1635
rect 200 1585 250 1615
rect 200 1565 215 1585
rect 235 1565 250 1585
rect 200 1535 250 1565
rect 200 1515 215 1535
rect 235 1515 250 1535
rect 200 1485 250 1515
rect 200 1465 215 1485
rect 235 1465 250 1485
rect 200 1435 250 1465
rect 200 1415 215 1435
rect 235 1415 250 1435
rect 200 1385 250 1415
rect 200 1365 215 1385
rect 235 1365 250 1385
rect 200 1335 250 1365
rect 200 1315 215 1335
rect 235 1315 250 1335
rect 200 1285 250 1315
rect 200 1265 215 1285
rect 235 1265 250 1285
rect 200 1235 250 1265
rect 200 1215 215 1235
rect 235 1215 250 1235
rect 200 1185 250 1215
rect 200 1165 215 1185
rect 235 1165 250 1185
rect 200 1150 250 1165
<< pdiff >>
rect 0 3585 50 3600
rect 0 3565 15 3585
rect 35 3565 50 3585
rect 0 3535 50 3565
rect 0 3515 15 3535
rect 35 3515 50 3535
rect 0 3485 50 3515
rect 0 3465 15 3485
rect 35 3465 50 3485
rect 0 3435 50 3465
rect 0 3415 15 3435
rect 35 3415 50 3435
rect 0 3385 50 3415
rect 0 3365 15 3385
rect 35 3365 50 3385
rect 0 3335 50 3365
rect 0 3315 15 3335
rect 35 3315 50 3335
rect 0 3285 50 3315
rect 0 3265 15 3285
rect 35 3265 50 3285
rect 0 3235 50 3265
rect 0 3215 15 3235
rect 35 3215 50 3235
rect 0 3185 50 3215
rect 0 3165 15 3185
rect 35 3165 50 3185
rect 0 3135 50 3165
rect 0 3115 15 3135
rect 35 3115 50 3135
rect 0 3100 50 3115
rect 100 3585 150 3600
rect 100 3565 115 3585
rect 135 3565 150 3585
rect 100 3535 150 3565
rect 100 3515 115 3535
rect 135 3515 150 3535
rect 100 3485 150 3515
rect 100 3465 115 3485
rect 135 3465 150 3485
rect 100 3435 150 3465
rect 100 3415 115 3435
rect 135 3415 150 3435
rect 100 3385 150 3415
rect 100 3365 115 3385
rect 135 3365 150 3385
rect 100 3335 150 3365
rect 100 3315 115 3335
rect 135 3315 150 3335
rect 100 3285 150 3315
rect 100 3265 115 3285
rect 135 3265 150 3285
rect 100 3235 150 3265
rect 100 3215 115 3235
rect 135 3215 150 3235
rect 100 3185 150 3215
rect 100 3165 115 3185
rect 135 3165 150 3185
rect 100 3135 150 3165
rect 100 3115 115 3135
rect 135 3115 150 3135
rect 100 3100 150 3115
rect 200 3585 250 3600
rect 200 3565 215 3585
rect 235 3565 250 3585
rect 200 3535 250 3565
rect 200 3515 215 3535
rect 235 3515 250 3535
rect 200 3485 250 3515
rect 200 3465 215 3485
rect 235 3465 250 3485
rect 200 3435 250 3465
rect 200 3415 215 3435
rect 235 3415 250 3435
rect 200 3385 250 3415
rect 200 3365 215 3385
rect 235 3365 250 3385
rect 200 3335 250 3365
rect 200 3315 215 3335
rect 235 3315 250 3335
rect 200 3285 250 3315
rect 200 3265 215 3285
rect 235 3265 250 3285
rect 200 3235 250 3265
rect 200 3215 215 3235
rect 235 3215 250 3235
rect 200 3185 250 3215
rect 200 3165 215 3185
rect 235 3165 250 3185
rect 200 3135 250 3165
rect 200 3115 215 3135
rect 235 3115 250 3135
rect 200 3100 250 3115
rect 0 735 50 750
rect 0 715 15 735
rect 35 715 50 735
rect 0 685 50 715
rect 0 665 15 685
rect 35 665 50 685
rect 0 635 50 665
rect 0 615 15 635
rect 35 615 50 635
rect 0 585 50 615
rect 0 565 15 585
rect 35 565 50 585
rect 0 535 50 565
rect 0 515 15 535
rect 35 515 50 535
rect 0 485 50 515
rect 0 465 15 485
rect 35 465 50 485
rect 0 435 50 465
rect 0 415 15 435
rect 35 415 50 435
rect 0 385 50 415
rect 0 365 15 385
rect 35 365 50 385
rect 0 335 50 365
rect 0 315 15 335
rect 35 315 50 335
rect 0 285 50 315
rect 0 265 15 285
rect 35 265 50 285
rect 0 250 50 265
rect 100 735 150 750
rect 100 715 115 735
rect 135 715 150 735
rect 100 685 150 715
rect 100 665 115 685
rect 135 665 150 685
rect 100 635 150 665
rect 100 615 115 635
rect 135 615 150 635
rect 100 585 150 615
rect 100 565 115 585
rect 135 565 150 585
rect 100 535 150 565
rect 100 515 115 535
rect 135 515 150 535
rect 100 485 150 515
rect 100 465 115 485
rect 135 465 150 485
rect 100 435 150 465
rect 100 415 115 435
rect 135 415 150 435
rect 100 385 150 415
rect 100 365 115 385
rect 135 365 150 385
rect 100 335 150 365
rect 100 315 115 335
rect 135 315 150 335
rect 100 285 150 315
rect 100 265 115 285
rect 135 265 150 285
rect 100 250 150 265
rect 200 735 250 750
rect 200 715 215 735
rect 235 715 250 735
rect 200 685 250 715
rect 200 665 215 685
rect 235 665 250 685
rect 200 635 250 665
rect 200 615 215 635
rect 235 615 250 635
rect 200 585 250 615
rect 200 565 215 585
rect 235 565 250 585
rect 200 535 250 565
rect 200 515 215 535
rect 235 515 250 535
rect 200 485 250 515
rect 200 465 215 485
rect 235 465 250 485
rect 200 435 250 465
rect 200 415 215 435
rect 235 415 250 435
rect 200 385 250 415
rect 200 365 215 385
rect 235 365 250 385
rect 200 335 250 365
rect 200 315 215 335
rect 235 315 250 335
rect 200 285 250 315
rect 200 265 215 285
rect 235 265 250 285
rect 200 250 250 265
<< ndiffc >>
rect 15 2665 35 2685
rect 15 2615 35 2635
rect 15 2565 35 2585
rect 15 2515 35 2535
rect 15 2465 35 2485
rect 15 2415 35 2435
rect 15 2365 35 2385
rect 15 2315 35 2335
rect 15 2265 35 2285
rect 15 2215 35 2235
rect 15 2165 35 2185
rect 15 2115 35 2135
rect 15 2065 35 2085
rect 15 2015 35 2035
rect 115 2665 135 2685
rect 115 2615 135 2635
rect 115 2565 135 2585
rect 115 2515 135 2535
rect 115 2465 135 2485
rect 115 2415 135 2435
rect 115 2365 135 2385
rect 115 2315 135 2335
rect 115 2265 135 2285
rect 115 2215 135 2235
rect 115 2165 135 2185
rect 115 2115 135 2135
rect 115 2065 135 2085
rect 115 2015 135 2035
rect 215 2665 235 2685
rect 215 2615 235 2635
rect 215 2565 235 2585
rect 215 2515 235 2535
rect 215 2465 235 2485
rect 215 2415 235 2435
rect 215 2365 235 2385
rect 215 2315 235 2335
rect 215 2265 235 2285
rect 215 2215 235 2235
rect 215 2165 235 2185
rect 215 2115 235 2135
rect 215 2065 235 2085
rect 215 2015 235 2035
rect 15 1815 35 1835
rect 15 1765 35 1785
rect 15 1715 35 1735
rect 15 1665 35 1685
rect 15 1615 35 1635
rect 15 1565 35 1585
rect 15 1515 35 1535
rect 15 1465 35 1485
rect 15 1415 35 1435
rect 15 1365 35 1385
rect 15 1315 35 1335
rect 15 1265 35 1285
rect 15 1215 35 1235
rect 15 1165 35 1185
rect 115 1815 135 1835
rect 115 1765 135 1785
rect 115 1715 135 1735
rect 115 1665 135 1685
rect 115 1615 135 1635
rect 115 1565 135 1585
rect 115 1515 135 1535
rect 115 1465 135 1485
rect 115 1415 135 1435
rect 115 1365 135 1385
rect 115 1315 135 1335
rect 115 1265 135 1285
rect 115 1215 135 1235
rect 115 1165 135 1185
rect 215 1815 235 1835
rect 215 1765 235 1785
rect 215 1715 235 1735
rect 215 1665 235 1685
rect 215 1615 235 1635
rect 215 1565 235 1585
rect 215 1515 235 1535
rect 215 1465 235 1485
rect 215 1415 235 1435
rect 215 1365 235 1385
rect 215 1315 235 1335
rect 215 1265 235 1285
rect 215 1215 235 1235
rect 215 1165 235 1185
<< pdiffc >>
rect 15 3565 35 3585
rect 15 3515 35 3535
rect 15 3465 35 3485
rect 15 3415 35 3435
rect 15 3365 35 3385
rect 15 3315 35 3335
rect 15 3265 35 3285
rect 15 3215 35 3235
rect 15 3165 35 3185
rect 15 3115 35 3135
rect 115 3565 135 3585
rect 115 3515 135 3535
rect 115 3465 135 3485
rect 115 3415 135 3435
rect 115 3365 135 3385
rect 115 3315 135 3335
rect 115 3265 135 3285
rect 115 3215 135 3235
rect 115 3165 135 3185
rect 115 3115 135 3135
rect 215 3565 235 3585
rect 215 3515 235 3535
rect 215 3465 235 3485
rect 215 3415 235 3435
rect 215 3365 235 3385
rect 215 3315 235 3335
rect 215 3265 235 3285
rect 215 3215 235 3235
rect 215 3165 235 3185
rect 215 3115 235 3135
rect 15 715 35 735
rect 15 665 35 685
rect 15 615 35 635
rect 15 565 35 585
rect 15 515 35 535
rect 15 465 35 485
rect 15 415 35 435
rect 15 365 35 385
rect 15 315 35 335
rect 15 265 35 285
rect 115 715 135 735
rect 115 665 135 685
rect 115 615 135 635
rect 115 565 135 585
rect 115 515 135 535
rect 115 465 135 485
rect 115 415 135 435
rect 115 365 135 385
rect 115 315 135 335
rect 115 265 135 285
rect 215 715 235 735
rect 215 665 235 685
rect 215 615 235 635
rect 215 565 235 585
rect 215 515 235 535
rect 215 465 235 485
rect 215 415 235 435
rect 215 365 235 385
rect 215 315 235 335
rect 215 265 235 285
<< psubdiff >>
rect -50 3835 300 3850
rect -50 3815 -35 3835
rect -15 3815 15 3835
rect 35 3815 65 3835
rect 85 3815 115 3835
rect 135 3815 165 3835
rect 185 3815 215 3835
rect 235 3815 265 3835
rect 285 3815 300 3835
rect -50 3800 300 3815
rect 0 2785 250 2800
rect 0 2765 15 2785
rect 35 2765 65 2785
rect 85 2765 115 2785
rect 135 2765 165 2785
rect 185 2765 215 2785
rect 235 2765 250 2785
rect 0 2750 250 2765
rect 0 1085 250 1100
rect 0 1065 15 1085
rect 35 1065 65 1085
rect 85 1065 115 1085
rect 135 1065 165 1085
rect 185 1065 215 1085
rect 235 1065 250 1085
rect 0 1050 250 1065
rect -50 35 300 50
rect -50 15 -35 35
rect -15 15 15 35
rect 35 15 65 35
rect 85 15 115 35
rect 135 15 165 35
rect 185 15 215 35
rect 235 15 265 35
rect 285 15 300 35
rect -50 0 300 15
<< nsubdiff >>
rect 0 3685 250 3700
rect 0 3665 15 3685
rect 35 3665 65 3685
rect 85 3665 115 3685
rect 135 3665 165 3685
rect 185 3665 215 3685
rect 235 3665 250 3685
rect 0 3650 250 3665
rect 0 2935 250 2950
rect 0 2915 15 2935
rect 35 2915 65 2935
rect 85 2915 115 2935
rect 135 2915 165 2935
rect 185 2915 215 2935
rect 235 2915 250 2935
rect 0 2900 250 2915
rect 0 935 250 950
rect 0 915 15 935
rect 35 915 65 935
rect 85 915 115 935
rect 135 915 165 935
rect 185 915 215 935
rect 235 915 250 935
rect 0 900 250 915
rect 0 185 250 200
rect 0 165 15 185
rect 35 165 65 185
rect 85 165 115 185
rect 135 165 165 185
rect 185 165 215 185
rect 235 165 250 185
rect 0 150 250 165
<< psubdiffcont >>
rect -35 3815 -15 3835
rect 15 3815 35 3835
rect 65 3815 85 3835
rect 115 3815 135 3835
rect 165 3815 185 3835
rect 215 3815 235 3835
rect 265 3815 285 3835
rect 15 2765 35 2785
rect 65 2765 85 2785
rect 115 2765 135 2785
rect 165 2765 185 2785
rect 215 2765 235 2785
rect 15 1065 35 1085
rect 65 1065 85 1085
rect 115 1065 135 1085
rect 165 1065 185 1085
rect 215 1065 235 1085
rect -35 15 -15 35
rect 15 15 35 35
rect 65 15 85 35
rect 115 15 135 35
rect 165 15 185 35
rect 215 15 235 35
rect 265 15 285 35
<< nsubdiffcont >>
rect 15 3665 35 3685
rect 65 3665 85 3685
rect 115 3665 135 3685
rect 165 3665 185 3685
rect 215 3665 235 3685
rect 15 2915 35 2935
rect 65 2915 85 2935
rect 115 2915 135 2935
rect 165 2915 185 2935
rect 215 2915 235 2935
rect 15 915 35 935
rect 65 915 85 935
rect 115 915 135 935
rect 165 915 185 935
rect 215 915 235 935
rect 15 165 35 185
rect 65 165 85 185
rect 115 165 135 185
rect 165 165 185 185
rect 215 165 235 185
<< poly >>
rect 50 3600 100 3615
rect 150 3600 200 3615
rect 50 3050 100 3100
rect 150 3050 200 3100
rect 50 3035 200 3050
rect 50 3015 65 3035
rect 85 3015 115 3035
rect 135 3015 165 3035
rect 185 3015 200 3035
rect 50 3000 200 3015
rect 50 2700 100 2715
rect 150 2700 200 2715
rect 50 1950 100 2000
rect 150 1950 200 2000
rect 50 1935 200 1950
rect 50 1915 65 1935
rect 85 1915 115 1935
rect 135 1915 165 1935
rect 185 1915 200 1935
rect 50 1900 200 1915
rect 50 1850 100 1900
rect 150 1850 200 1900
rect 50 1135 100 1150
rect 150 1135 200 1150
rect 50 835 200 850
rect 50 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 200 835
rect 50 800 200 815
rect 50 750 100 800
rect 150 750 200 800
rect 50 235 100 250
rect 150 235 200 250
<< polycont >>
rect 65 3015 85 3035
rect 115 3015 135 3035
rect 165 3015 185 3035
rect 65 1915 85 1935
rect 115 1915 135 1935
rect 165 1915 185 1935
rect 65 815 85 835
rect 115 815 135 835
rect 165 815 185 835
<< locali >>
rect -50 3835 300 3850
rect -50 3815 -35 3835
rect -15 3815 15 3835
rect 35 3815 65 3835
rect 85 3815 115 3835
rect 135 3815 165 3835
rect 185 3815 215 3835
rect 235 3815 265 3835
rect 285 3815 300 3835
rect -50 3800 300 3815
rect 0 3685 250 3700
rect 0 3665 15 3685
rect 35 3665 65 3685
rect 85 3665 115 3685
rect 135 3665 165 3685
rect 185 3665 215 3685
rect 235 3665 250 3685
rect 0 3650 250 3665
rect 0 3585 50 3600
rect 0 3565 15 3585
rect 35 3565 50 3585
rect 0 3535 50 3565
rect 0 3515 15 3535
rect 35 3515 50 3535
rect 0 3485 50 3515
rect 0 3465 15 3485
rect 35 3465 50 3485
rect 0 3435 50 3465
rect 0 3415 15 3435
rect 35 3415 50 3435
rect 0 3385 50 3415
rect 0 3365 15 3385
rect 35 3365 50 3385
rect 0 3335 50 3365
rect 0 3315 15 3335
rect 35 3315 50 3335
rect 0 3285 50 3315
rect 0 3265 15 3285
rect 35 3265 50 3285
rect 0 3235 50 3265
rect 0 3215 15 3235
rect 35 3215 50 3235
rect 0 3185 50 3215
rect 0 3165 15 3185
rect 35 3165 50 3185
rect 0 3135 50 3165
rect 0 3115 15 3135
rect 35 3115 50 3135
rect 0 3100 50 3115
rect 100 3585 150 3600
rect 100 3565 115 3585
rect 135 3565 150 3585
rect 100 3535 150 3565
rect 100 3515 115 3535
rect 135 3515 150 3535
rect 100 3485 150 3515
rect 100 3465 115 3485
rect 135 3465 150 3485
rect 100 3435 150 3465
rect 100 3415 115 3435
rect 135 3415 150 3435
rect 100 3385 150 3415
rect 100 3365 115 3385
rect 135 3365 150 3385
rect 100 3335 150 3365
rect 100 3315 115 3335
rect 135 3315 150 3335
rect 100 3285 150 3315
rect 100 3265 115 3285
rect 135 3265 150 3285
rect 100 3235 150 3265
rect 100 3215 115 3235
rect 135 3215 150 3235
rect 100 3185 150 3215
rect 100 3165 115 3185
rect 135 3165 150 3185
rect 100 3135 150 3165
rect 100 3115 115 3135
rect 135 3115 150 3135
rect 100 3100 150 3115
rect 200 3585 250 3600
rect 200 3565 215 3585
rect 235 3565 250 3585
rect 200 3535 250 3565
rect 200 3515 215 3535
rect 235 3515 250 3535
rect 200 3485 250 3515
rect 200 3465 215 3485
rect 235 3465 250 3485
rect 200 3435 250 3465
rect 200 3415 215 3435
rect 235 3415 250 3435
rect 200 3385 250 3415
rect 200 3365 215 3385
rect 235 3365 250 3385
rect 200 3335 250 3365
rect 200 3315 215 3335
rect 235 3315 250 3335
rect 200 3285 250 3315
rect 200 3265 215 3285
rect 235 3265 250 3285
rect 200 3235 250 3265
rect 200 3215 215 3235
rect 235 3215 250 3235
rect 200 3185 250 3215
rect 200 3165 215 3185
rect 235 3165 250 3185
rect 200 3135 250 3165
rect 200 3115 215 3135
rect 235 3115 250 3135
rect 200 3100 250 3115
rect 50 3035 200 3050
rect 50 3015 65 3035
rect 85 3015 115 3035
rect 135 3015 165 3035
rect 185 3015 200 3035
rect 50 3000 200 3015
rect 0 2935 250 2950
rect 0 2915 15 2935
rect 35 2915 65 2935
rect 85 2915 115 2935
rect 135 2915 165 2935
rect 185 2915 215 2935
rect 235 2915 250 2935
rect 0 2900 250 2915
rect 0 2785 250 2800
rect 0 2765 15 2785
rect 35 2765 65 2785
rect 85 2765 115 2785
rect 135 2765 165 2785
rect 185 2765 215 2785
rect 235 2765 250 2785
rect 0 2750 250 2765
rect 0 2685 50 2700
rect 0 2665 15 2685
rect 35 2665 50 2685
rect 0 2635 50 2665
rect 0 2615 15 2635
rect 35 2615 50 2635
rect 0 2585 50 2615
rect 0 2565 15 2585
rect 35 2565 50 2585
rect 0 2535 50 2565
rect 0 2515 15 2535
rect 35 2515 50 2535
rect 0 2485 50 2515
rect 0 2465 15 2485
rect 35 2465 50 2485
rect 0 2435 50 2465
rect 0 2415 15 2435
rect 35 2415 50 2435
rect 0 2385 50 2415
rect 0 2365 15 2385
rect 35 2365 50 2385
rect 0 2335 50 2365
rect 0 2315 15 2335
rect 35 2315 50 2335
rect 0 2285 50 2315
rect 0 2265 15 2285
rect 35 2265 50 2285
rect 0 2235 50 2265
rect 0 2215 15 2235
rect 35 2215 50 2235
rect 0 2185 50 2215
rect 0 2165 15 2185
rect 35 2165 50 2185
rect 0 2135 50 2165
rect 0 2115 15 2135
rect 35 2115 50 2135
rect 0 2085 50 2115
rect 0 2065 15 2085
rect 35 2065 50 2085
rect 0 2035 50 2065
rect 0 2015 15 2035
rect 35 2015 50 2035
rect 0 2000 50 2015
rect 100 2685 150 2700
rect 100 2665 115 2685
rect 135 2665 150 2685
rect 100 2635 150 2665
rect 100 2615 115 2635
rect 135 2615 150 2635
rect 100 2585 150 2615
rect 100 2565 115 2585
rect 135 2565 150 2585
rect 100 2535 150 2565
rect 100 2515 115 2535
rect 135 2515 150 2535
rect 100 2485 150 2515
rect 100 2465 115 2485
rect 135 2465 150 2485
rect 100 2435 150 2465
rect 100 2415 115 2435
rect 135 2415 150 2435
rect 100 2385 150 2415
rect 100 2365 115 2385
rect 135 2365 150 2385
rect 100 2335 150 2365
rect 100 2315 115 2335
rect 135 2315 150 2335
rect 100 2285 150 2315
rect 100 2265 115 2285
rect 135 2265 150 2285
rect 100 2235 150 2265
rect 100 2215 115 2235
rect 135 2215 150 2235
rect 100 2185 150 2215
rect 100 2165 115 2185
rect 135 2165 150 2185
rect 100 2135 150 2165
rect 100 2115 115 2135
rect 135 2115 150 2135
rect 100 2085 150 2115
rect 100 2065 115 2085
rect 135 2065 150 2085
rect 100 2035 150 2065
rect 100 2015 115 2035
rect 135 2015 150 2035
rect 100 2000 150 2015
rect 200 2685 250 2700
rect 200 2665 215 2685
rect 235 2665 250 2685
rect 200 2635 250 2665
rect 200 2615 215 2635
rect 235 2615 250 2635
rect 200 2585 250 2615
rect 200 2565 215 2585
rect 235 2565 250 2585
rect 200 2535 250 2565
rect 200 2515 215 2535
rect 235 2515 250 2535
rect 200 2485 250 2515
rect 200 2465 215 2485
rect 235 2465 250 2485
rect 200 2435 250 2465
rect 200 2415 215 2435
rect 235 2415 250 2435
rect 200 2385 250 2415
rect 200 2365 215 2385
rect 235 2365 250 2385
rect 200 2335 250 2365
rect 200 2315 215 2335
rect 235 2315 250 2335
rect 200 2285 250 2315
rect 200 2265 215 2285
rect 235 2265 250 2285
rect 200 2235 250 2265
rect 200 2215 215 2235
rect 235 2215 250 2235
rect 200 2185 250 2215
rect 200 2165 215 2185
rect 235 2165 250 2185
rect 200 2135 250 2165
rect 200 2115 215 2135
rect 235 2115 250 2135
rect 200 2085 250 2115
rect 200 2065 215 2085
rect 235 2065 250 2085
rect 200 2035 250 2065
rect 200 2015 215 2035
rect 235 2015 250 2035
rect 200 2000 250 2015
rect 50 1935 200 1950
rect 50 1915 65 1935
rect 85 1915 115 1935
rect 135 1915 165 1935
rect 185 1915 200 1935
rect 50 1900 200 1915
rect 0 1835 50 1850
rect 0 1815 15 1835
rect 35 1815 50 1835
rect 0 1785 50 1815
rect 0 1765 15 1785
rect 35 1765 50 1785
rect 0 1735 50 1765
rect 0 1715 15 1735
rect 35 1715 50 1735
rect 0 1685 50 1715
rect 0 1665 15 1685
rect 35 1665 50 1685
rect 0 1635 50 1665
rect 0 1615 15 1635
rect 35 1615 50 1635
rect 0 1585 50 1615
rect 0 1565 15 1585
rect 35 1565 50 1585
rect 0 1535 50 1565
rect 0 1515 15 1535
rect 35 1515 50 1535
rect 0 1485 50 1515
rect 0 1465 15 1485
rect 35 1465 50 1485
rect 0 1435 50 1465
rect 0 1415 15 1435
rect 35 1415 50 1435
rect 0 1385 50 1415
rect 0 1365 15 1385
rect 35 1365 50 1385
rect 0 1335 50 1365
rect 0 1315 15 1335
rect 35 1315 50 1335
rect 0 1285 50 1315
rect 0 1265 15 1285
rect 35 1265 50 1285
rect 0 1235 50 1265
rect 0 1215 15 1235
rect 35 1215 50 1235
rect 0 1185 50 1215
rect 0 1165 15 1185
rect 35 1165 50 1185
rect 0 1150 50 1165
rect 100 1835 150 1850
rect 100 1815 115 1835
rect 135 1815 150 1835
rect 100 1785 150 1815
rect 100 1765 115 1785
rect 135 1765 150 1785
rect 100 1735 150 1765
rect 100 1715 115 1735
rect 135 1715 150 1735
rect 100 1685 150 1715
rect 100 1665 115 1685
rect 135 1665 150 1685
rect 100 1635 150 1665
rect 100 1615 115 1635
rect 135 1615 150 1635
rect 100 1585 150 1615
rect 100 1565 115 1585
rect 135 1565 150 1585
rect 100 1535 150 1565
rect 100 1515 115 1535
rect 135 1515 150 1535
rect 100 1485 150 1515
rect 100 1465 115 1485
rect 135 1465 150 1485
rect 100 1435 150 1465
rect 100 1415 115 1435
rect 135 1415 150 1435
rect 100 1385 150 1415
rect 100 1365 115 1385
rect 135 1365 150 1385
rect 100 1335 150 1365
rect 100 1315 115 1335
rect 135 1315 150 1335
rect 100 1285 150 1315
rect 100 1265 115 1285
rect 135 1265 150 1285
rect 100 1235 150 1265
rect 100 1215 115 1235
rect 135 1215 150 1235
rect 100 1185 150 1215
rect 100 1165 115 1185
rect 135 1165 150 1185
rect 100 1150 150 1165
rect 200 1835 250 1850
rect 200 1815 215 1835
rect 235 1815 250 1835
rect 200 1785 250 1815
rect 200 1765 215 1785
rect 235 1765 250 1785
rect 200 1735 250 1765
rect 200 1715 215 1735
rect 235 1715 250 1735
rect 200 1685 250 1715
rect 200 1665 215 1685
rect 235 1665 250 1685
rect 200 1635 250 1665
rect 200 1615 215 1635
rect 235 1615 250 1635
rect 200 1585 250 1615
rect 200 1565 215 1585
rect 235 1565 250 1585
rect 200 1535 250 1565
rect 200 1515 215 1535
rect 235 1515 250 1535
rect 200 1485 250 1515
rect 200 1465 215 1485
rect 235 1465 250 1485
rect 200 1435 250 1465
rect 200 1415 215 1435
rect 235 1415 250 1435
rect 200 1385 250 1415
rect 200 1365 215 1385
rect 235 1365 250 1385
rect 200 1335 250 1365
rect 200 1315 215 1335
rect 235 1315 250 1335
rect 200 1285 250 1315
rect 200 1265 215 1285
rect 235 1265 250 1285
rect 200 1235 250 1265
rect 200 1215 215 1235
rect 235 1215 250 1235
rect 200 1185 250 1215
rect 200 1165 215 1185
rect 235 1165 250 1185
rect 200 1150 250 1165
rect 0 1085 250 1100
rect 0 1065 15 1085
rect 35 1065 65 1085
rect 85 1065 115 1085
rect 135 1065 165 1085
rect 185 1065 215 1085
rect 235 1065 250 1085
rect 0 1050 250 1065
rect 0 935 250 950
rect 0 915 15 935
rect 35 915 65 935
rect 85 915 115 935
rect 135 915 165 935
rect 185 915 215 935
rect 235 915 250 935
rect 0 900 250 915
rect 50 835 200 850
rect 50 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 200 835
rect 50 800 200 815
rect 0 735 50 750
rect 0 715 15 735
rect 35 715 50 735
rect 0 685 50 715
rect 0 665 15 685
rect 35 665 50 685
rect 0 635 50 665
rect 0 615 15 635
rect 35 615 50 635
rect 0 585 50 615
rect 0 565 15 585
rect 35 565 50 585
rect 0 535 50 565
rect 0 515 15 535
rect 35 515 50 535
rect 0 485 50 515
rect 0 465 15 485
rect 35 465 50 485
rect 0 435 50 465
rect 0 415 15 435
rect 35 415 50 435
rect 0 385 50 415
rect 0 365 15 385
rect 35 365 50 385
rect 0 335 50 365
rect 0 315 15 335
rect 35 315 50 335
rect 0 285 50 315
rect 0 265 15 285
rect 35 265 50 285
rect 0 250 50 265
rect 100 735 150 750
rect 100 715 115 735
rect 135 715 150 735
rect 100 685 150 715
rect 100 665 115 685
rect 135 665 150 685
rect 100 635 150 665
rect 100 615 115 635
rect 135 615 150 635
rect 100 585 150 615
rect 100 565 115 585
rect 135 565 150 585
rect 100 535 150 565
rect 100 515 115 535
rect 135 515 150 535
rect 100 485 150 515
rect 100 465 115 485
rect 135 465 150 485
rect 100 435 150 465
rect 100 415 115 435
rect 135 415 150 435
rect 100 385 150 415
rect 100 365 115 385
rect 135 365 150 385
rect 100 335 150 365
rect 100 315 115 335
rect 135 315 150 335
rect 100 285 150 315
rect 100 265 115 285
rect 135 265 150 285
rect 100 250 150 265
rect 200 735 250 750
rect 200 715 215 735
rect 235 715 250 735
rect 200 685 250 715
rect 200 665 215 685
rect 235 665 250 685
rect 200 635 250 665
rect 200 615 215 635
rect 235 615 250 635
rect 200 585 250 615
rect 200 565 215 585
rect 235 565 250 585
rect 200 535 250 565
rect 200 515 215 535
rect 235 515 250 535
rect 200 485 250 515
rect 200 465 215 485
rect 235 465 250 485
rect 200 435 250 465
rect 200 415 215 435
rect 235 415 250 435
rect 200 385 250 415
rect 200 365 215 385
rect 235 365 250 385
rect 200 335 250 365
rect 200 315 215 335
rect 235 315 250 335
rect 200 285 250 315
rect 200 265 215 285
rect 235 265 250 285
rect 200 250 250 265
rect 0 185 250 200
rect 0 165 15 185
rect 35 165 65 185
rect 85 165 115 185
rect 135 165 165 185
rect 185 165 215 185
rect 235 165 250 185
rect 0 150 250 165
rect -50 35 300 50
rect -50 15 -35 35
rect -15 15 15 35
rect 35 15 65 35
rect 85 15 115 35
rect 135 15 165 35
rect 185 15 215 35
rect 235 15 265 35
rect 285 15 300 35
rect -50 0 300 15
<< viali >>
rect 15 3565 35 3585
rect 15 3515 35 3535
rect 15 3465 35 3485
rect 15 3415 35 3435
rect 15 3365 35 3385
rect 15 3315 35 3335
rect 15 3265 35 3285
rect 15 3215 35 3235
rect 15 3165 35 3185
rect 15 3115 35 3135
rect 115 3565 135 3585
rect 115 3515 135 3535
rect 115 3465 135 3485
rect 115 3415 135 3435
rect 115 3365 135 3385
rect 115 3315 135 3335
rect 115 3265 135 3285
rect 115 3215 135 3235
rect 115 3165 135 3185
rect 115 3115 135 3135
rect 215 3565 235 3585
rect 215 3515 235 3535
rect 215 3465 235 3485
rect 215 3415 235 3435
rect 215 3365 235 3385
rect 215 3315 235 3335
rect 215 3265 235 3285
rect 215 3215 235 3235
rect 115 3015 135 3035
rect 15 2665 35 2685
rect 15 2615 35 2635
rect 15 2565 35 2585
rect 15 2515 35 2535
rect 15 2465 35 2485
rect 15 2415 35 2435
rect 15 2365 35 2385
rect 15 2315 35 2335
rect 15 2265 35 2285
rect 15 2215 35 2235
rect 15 2165 35 2185
rect 15 2115 35 2135
rect 15 2065 35 2085
rect 15 2015 35 2035
rect 115 2665 135 2685
rect 115 2615 135 2635
rect 115 2565 135 2585
rect 115 2515 135 2535
rect 115 2465 135 2485
rect 115 2415 135 2435
rect 115 2365 135 2385
rect 115 2315 135 2335
rect 115 2265 135 2285
rect 115 2215 135 2235
rect 115 2165 135 2185
rect 115 2115 135 2135
rect 115 2065 135 2085
rect 115 2015 135 2035
rect 215 2665 235 2685
rect 215 2615 235 2635
rect 215 2565 235 2585
rect 215 2515 235 2535
rect 215 2465 235 2485
rect 215 2415 235 2435
rect 215 2365 235 2385
rect 215 2315 235 2335
rect 215 2265 235 2285
rect 215 2215 235 2235
rect 215 2165 235 2185
rect 215 2115 235 2135
rect 215 2065 235 2085
rect 215 2015 235 2035
rect 115 1915 135 1935
rect 15 1815 35 1835
rect 15 1765 35 1785
rect 15 1715 35 1735
rect 15 1665 35 1685
rect 15 1615 35 1635
rect 15 1565 35 1585
rect 15 1515 35 1535
rect 15 1465 35 1485
rect 15 1415 35 1435
rect 15 1365 35 1385
rect 15 1315 35 1335
rect 15 1265 35 1285
rect 15 1215 35 1235
rect 15 1165 35 1185
rect 115 1815 135 1835
rect 115 1765 135 1785
rect 115 1715 135 1735
rect 115 1665 135 1685
rect 115 1615 135 1635
rect 115 1565 135 1585
rect 115 1515 135 1535
rect 115 1465 135 1485
rect 115 1415 135 1435
rect 115 1365 135 1385
rect 115 1315 135 1335
rect 115 1265 135 1285
rect 115 1215 135 1235
rect 115 1165 135 1185
rect 215 1815 235 1835
rect 215 1765 235 1785
rect 215 1715 235 1735
rect 215 1665 235 1685
rect 215 1615 235 1635
rect 215 1565 235 1585
rect 215 1515 235 1535
rect 215 1465 235 1485
rect 215 1415 235 1435
rect 215 1365 235 1385
rect 215 1315 235 1335
rect 215 1265 235 1285
rect 215 1215 235 1235
rect 215 1165 235 1185
rect 115 815 135 835
rect 15 715 35 735
rect 15 665 35 685
rect 15 615 35 635
rect 15 565 35 585
rect 15 515 35 535
rect 15 465 35 485
rect 15 415 35 435
rect 15 365 35 385
rect 15 315 35 335
rect 15 265 35 285
rect 115 715 135 735
rect 115 665 135 685
rect 115 615 135 635
rect 115 565 135 585
rect 115 515 135 535
rect 115 465 135 485
rect 115 415 135 435
rect 115 365 135 385
rect 115 315 135 335
rect 115 265 135 285
rect 215 615 235 635
rect 215 565 235 585
rect 215 515 235 535
rect 215 465 235 485
rect 215 415 235 435
rect 215 365 235 385
rect 215 315 235 335
rect 215 265 235 285
<< metal1 >>
rect 0 3740 50 3750
rect 0 3710 10 3740
rect 40 3710 50 3740
rect 0 3640 50 3710
rect 0 3610 10 3640
rect 40 3610 50 3640
rect 0 3585 50 3610
rect 200 3740 250 3750
rect 200 3710 210 3740
rect 240 3710 250 3740
rect 200 3640 250 3710
rect 200 3610 210 3640
rect 240 3610 250 3640
rect 0 3565 15 3585
rect 35 3565 50 3585
rect 0 3540 50 3565
rect 0 3510 10 3540
rect 40 3510 50 3540
rect 0 3485 50 3510
rect 0 3465 15 3485
rect 35 3465 50 3485
rect 0 3440 50 3465
rect 0 3410 10 3440
rect 40 3410 50 3440
rect 0 3385 50 3410
rect 0 3365 15 3385
rect 35 3365 50 3385
rect 0 3340 50 3365
rect 0 3310 10 3340
rect 40 3310 50 3340
rect 0 3285 50 3310
rect 0 3265 15 3285
rect 35 3265 50 3285
rect 0 3240 50 3265
rect 0 3210 10 3240
rect 40 3210 50 3240
rect 0 3185 50 3210
rect 0 3165 15 3185
rect 35 3165 50 3185
rect 0 3140 50 3165
rect 0 3110 10 3140
rect 40 3110 50 3140
rect 0 3100 50 3110
rect 100 3585 150 3600
rect 100 3565 115 3585
rect 135 3565 150 3585
rect 100 3535 150 3565
rect 100 3515 115 3535
rect 135 3515 150 3535
rect 100 3485 150 3515
rect 100 3465 115 3485
rect 135 3465 150 3485
rect 100 3435 150 3465
rect 100 3415 115 3435
rect 135 3415 150 3435
rect 100 3385 150 3415
rect 100 3365 115 3385
rect 135 3365 150 3385
rect 100 3335 150 3365
rect 100 3315 115 3335
rect 135 3315 150 3335
rect 100 3285 150 3315
rect 100 3265 115 3285
rect 135 3265 150 3285
rect 100 3235 150 3265
rect 100 3215 115 3235
rect 135 3215 150 3235
rect 100 3185 150 3215
rect 200 3585 250 3610
rect 200 3565 215 3585
rect 235 3565 250 3585
rect 200 3540 250 3565
rect 200 3510 210 3540
rect 240 3510 250 3540
rect 200 3485 250 3510
rect 200 3465 215 3485
rect 235 3465 250 3485
rect 200 3440 250 3465
rect 200 3410 210 3440
rect 240 3410 250 3440
rect 200 3385 250 3410
rect 200 3365 215 3385
rect 235 3365 250 3385
rect 200 3340 250 3365
rect 200 3310 210 3340
rect 240 3310 250 3340
rect 200 3285 250 3310
rect 200 3265 215 3285
rect 235 3265 250 3285
rect 200 3240 250 3265
rect 200 3210 210 3240
rect 240 3210 250 3240
rect 200 3200 250 3210
rect 100 3165 115 3185
rect 135 3165 150 3185
rect 100 3135 150 3165
rect 100 3115 115 3135
rect 135 3115 150 3135
rect 100 3040 150 3115
rect 200 3100 250 3150
rect 100 3010 110 3040
rect 140 3010 150 3040
rect 100 3000 150 3010
rect 0 2840 50 2850
rect 0 2810 10 2840
rect 40 2810 50 2840
rect 0 2685 50 2810
rect 200 2840 250 2850
rect 200 2810 210 2840
rect 240 2810 250 2840
rect 0 2665 15 2685
rect 35 2665 50 2685
rect 0 2635 50 2665
rect 0 2615 15 2635
rect 35 2615 50 2635
rect 0 2585 50 2615
rect 0 2565 15 2585
rect 35 2565 50 2585
rect 0 2535 50 2565
rect 0 2515 15 2535
rect 35 2515 50 2535
rect 0 2485 50 2515
rect 0 2465 15 2485
rect 35 2465 50 2485
rect 0 2440 50 2465
rect 0 2410 10 2440
rect 40 2410 50 2440
rect 0 2385 50 2410
rect 0 2365 15 2385
rect 35 2365 50 2385
rect 0 2340 50 2365
rect 0 2310 10 2340
rect 40 2310 50 2340
rect 0 2285 50 2310
rect 0 2265 15 2285
rect 35 2265 50 2285
rect 0 2240 50 2265
rect 0 2210 10 2240
rect 40 2210 50 2240
rect 0 2185 50 2210
rect 0 2165 15 2185
rect 35 2165 50 2185
rect 0 2140 50 2165
rect 0 2110 10 2140
rect 40 2110 50 2140
rect 0 2085 50 2110
rect 0 2065 15 2085
rect 35 2065 50 2085
rect 0 2040 50 2065
rect 0 2010 10 2040
rect 40 2010 50 2040
rect 0 1840 50 2010
rect 0 1810 10 1840
rect 40 1810 50 1840
rect 0 1785 50 1810
rect 0 1765 15 1785
rect 35 1765 50 1785
rect 0 1740 50 1765
rect 0 1710 10 1740
rect 40 1710 50 1740
rect 0 1685 50 1710
rect 0 1665 15 1685
rect 35 1665 50 1685
rect 0 1640 50 1665
rect 0 1610 10 1640
rect 40 1610 50 1640
rect 0 1585 50 1610
rect 0 1565 15 1585
rect 35 1565 50 1585
rect 0 1540 50 1565
rect 0 1510 10 1540
rect 40 1510 50 1540
rect 0 1485 50 1510
rect 0 1465 15 1485
rect 35 1465 50 1485
rect 0 1440 50 1465
rect 0 1410 10 1440
rect 40 1410 50 1440
rect 0 1385 50 1410
rect 0 1365 15 1385
rect 35 1365 50 1385
rect 0 1335 50 1365
rect 0 1315 15 1335
rect 35 1315 50 1335
rect 0 1285 50 1315
rect 0 1265 15 1285
rect 35 1265 50 1285
rect 0 1235 50 1265
rect 0 1215 15 1235
rect 35 1215 50 1235
rect 0 1185 50 1215
rect 0 1165 15 1185
rect 35 1165 50 1185
rect 0 1040 50 1165
rect 100 2685 150 2700
rect 100 2665 115 2685
rect 135 2665 150 2685
rect 100 2635 150 2665
rect 100 2615 115 2635
rect 135 2615 150 2635
rect 100 2585 150 2615
rect 100 2565 115 2585
rect 135 2565 150 2585
rect 100 2535 150 2565
rect 100 2515 115 2535
rect 135 2515 150 2535
rect 100 2485 150 2515
rect 100 2465 115 2485
rect 135 2465 150 2485
rect 100 2435 150 2465
rect 100 2415 115 2435
rect 135 2415 150 2435
rect 100 2385 150 2415
rect 100 2365 115 2385
rect 135 2365 150 2385
rect 100 2335 150 2365
rect 100 2315 115 2335
rect 135 2315 150 2335
rect 100 2285 150 2315
rect 100 2265 115 2285
rect 135 2265 150 2285
rect 100 2235 150 2265
rect 100 2215 115 2235
rect 135 2215 150 2235
rect 100 2185 150 2215
rect 100 2165 115 2185
rect 135 2165 150 2185
rect 100 2135 150 2165
rect 100 2115 115 2135
rect 135 2115 150 2135
rect 100 2085 150 2115
rect 100 2065 115 2085
rect 135 2065 150 2085
rect 100 2035 150 2065
rect 100 2015 115 2035
rect 135 2015 150 2035
rect 100 1940 150 2015
rect 100 1910 110 1940
rect 140 1910 150 1940
rect 100 1835 150 1910
rect 100 1815 115 1835
rect 135 1815 150 1835
rect 100 1785 150 1815
rect 100 1765 115 1785
rect 135 1765 150 1785
rect 100 1735 150 1765
rect 100 1715 115 1735
rect 135 1715 150 1735
rect 100 1685 150 1715
rect 100 1665 115 1685
rect 135 1665 150 1685
rect 100 1635 150 1665
rect 100 1615 115 1635
rect 135 1615 150 1635
rect 100 1585 150 1615
rect 100 1565 115 1585
rect 135 1565 150 1585
rect 100 1535 150 1565
rect 100 1515 115 1535
rect 135 1515 150 1535
rect 100 1485 150 1515
rect 100 1465 115 1485
rect 135 1465 150 1485
rect 100 1435 150 1465
rect 100 1415 115 1435
rect 135 1415 150 1435
rect 100 1385 150 1415
rect 100 1365 115 1385
rect 135 1365 150 1385
rect 100 1335 150 1365
rect 100 1315 115 1335
rect 135 1315 150 1335
rect 100 1285 150 1315
rect 100 1265 115 1285
rect 135 1265 150 1285
rect 100 1235 150 1265
rect 100 1215 115 1235
rect 135 1215 150 1235
rect 100 1185 150 1215
rect 100 1165 115 1185
rect 135 1165 150 1185
rect 100 1150 150 1165
rect 200 2685 250 2810
rect 200 2665 215 2685
rect 235 2665 250 2685
rect 200 2635 250 2665
rect 200 2615 215 2635
rect 235 2615 250 2635
rect 200 2585 250 2615
rect 200 2565 215 2585
rect 235 2565 250 2585
rect 200 2535 250 2565
rect 200 2515 215 2535
rect 235 2515 250 2535
rect 200 2485 250 2515
rect 200 2465 215 2485
rect 235 2465 250 2485
rect 200 2440 250 2465
rect 200 2410 210 2440
rect 240 2410 250 2440
rect 200 2385 250 2410
rect 200 2365 215 2385
rect 235 2365 250 2385
rect 200 2340 250 2365
rect 200 2310 210 2340
rect 240 2310 250 2340
rect 200 2285 250 2310
rect 200 2265 215 2285
rect 235 2265 250 2285
rect 200 2240 250 2265
rect 200 2210 210 2240
rect 240 2210 250 2240
rect 200 2185 250 2210
rect 200 2165 215 2185
rect 235 2165 250 2185
rect 200 2140 250 2165
rect 200 2110 210 2140
rect 240 2110 250 2140
rect 200 2085 250 2110
rect 200 2065 215 2085
rect 235 2065 250 2085
rect 200 2040 250 2065
rect 200 2010 210 2040
rect 240 2010 250 2040
rect 200 1840 250 2010
rect 200 1810 210 1840
rect 240 1810 250 1840
rect 200 1785 250 1810
rect 200 1765 215 1785
rect 235 1765 250 1785
rect 200 1740 250 1765
rect 200 1710 210 1740
rect 240 1710 250 1740
rect 200 1685 250 1710
rect 200 1665 215 1685
rect 235 1665 250 1685
rect 200 1640 250 1665
rect 200 1610 210 1640
rect 240 1610 250 1640
rect 200 1585 250 1610
rect 200 1565 215 1585
rect 235 1565 250 1585
rect 200 1540 250 1565
rect 200 1510 210 1540
rect 240 1510 250 1540
rect 200 1485 250 1510
rect 200 1465 215 1485
rect 235 1465 250 1485
rect 200 1440 250 1465
rect 200 1410 210 1440
rect 240 1410 250 1440
rect 200 1385 250 1410
rect 200 1365 215 1385
rect 235 1365 250 1385
rect 200 1335 250 1365
rect 200 1315 215 1335
rect 235 1315 250 1335
rect 200 1285 250 1315
rect 200 1265 215 1285
rect 235 1265 250 1285
rect 200 1235 250 1265
rect 200 1215 215 1235
rect 235 1215 250 1235
rect 200 1185 250 1215
rect 200 1165 215 1185
rect 235 1165 250 1185
rect 0 1010 10 1040
rect 40 1010 50 1040
rect 0 1000 50 1010
rect 200 1040 250 1165
rect 200 1010 210 1040
rect 240 1010 250 1040
rect 200 1000 250 1010
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 0 740 50 750
rect 0 710 10 740
rect 40 710 50 740
rect 0 685 50 710
rect 0 665 15 685
rect 35 665 50 685
rect 0 640 50 665
rect 0 610 10 640
rect 40 610 50 640
rect 0 585 50 610
rect 0 565 15 585
rect 35 565 50 585
rect 0 540 50 565
rect 0 510 10 540
rect 40 510 50 540
rect 0 485 50 510
rect 0 465 15 485
rect 35 465 50 485
rect 0 440 50 465
rect 0 410 10 440
rect 40 410 50 440
rect 0 385 50 410
rect 0 365 15 385
rect 35 365 50 385
rect 0 340 50 365
rect 0 310 10 340
rect 40 310 50 340
rect 0 285 50 310
rect 0 265 15 285
rect 35 265 50 285
rect 0 240 50 265
rect 100 735 150 810
rect 100 715 115 735
rect 135 715 150 735
rect 100 685 150 715
rect 200 700 250 750
rect 100 665 115 685
rect 135 665 150 685
rect 100 635 150 665
rect 100 615 115 635
rect 135 615 150 635
rect 100 585 150 615
rect 100 565 115 585
rect 135 565 150 585
rect 100 535 150 565
rect 100 515 115 535
rect 135 515 150 535
rect 100 485 150 515
rect 100 465 115 485
rect 135 465 150 485
rect 100 435 150 465
rect 100 415 115 435
rect 135 415 150 435
rect 100 385 150 415
rect 100 365 115 385
rect 135 365 150 385
rect 100 335 150 365
rect 100 315 115 335
rect 135 315 150 335
rect 100 285 150 315
rect 100 265 115 285
rect 135 265 150 285
rect 100 250 150 265
rect 200 640 250 650
rect 200 610 210 640
rect 240 610 250 640
rect 200 585 250 610
rect 200 565 215 585
rect 235 565 250 585
rect 200 540 250 565
rect 200 510 210 540
rect 240 510 250 540
rect 200 485 250 510
rect 200 465 215 485
rect 235 465 250 485
rect 200 440 250 465
rect 200 410 210 440
rect 240 410 250 440
rect 200 385 250 410
rect 200 365 215 385
rect 235 365 250 385
rect 200 340 250 365
rect 200 310 210 340
rect 240 310 250 340
rect 200 285 250 310
rect 200 265 215 285
rect 235 265 250 285
rect 0 210 10 240
rect 40 210 50 240
rect 0 140 50 210
rect 0 110 10 140
rect 40 110 50 140
rect 0 100 50 110
rect 200 240 250 265
rect 200 210 210 240
rect 240 210 250 240
rect 200 140 250 210
rect 200 110 210 140
rect 240 110 250 140
rect 200 100 250 110
<< via1 >>
rect 10 3710 40 3740
rect 10 3610 40 3640
rect 210 3710 240 3740
rect 210 3610 240 3640
rect 10 3535 40 3540
rect 10 3515 15 3535
rect 15 3515 35 3535
rect 35 3515 40 3535
rect 10 3510 40 3515
rect 10 3435 40 3440
rect 10 3415 15 3435
rect 15 3415 35 3435
rect 35 3415 40 3435
rect 10 3410 40 3415
rect 10 3335 40 3340
rect 10 3315 15 3335
rect 15 3315 35 3335
rect 35 3315 40 3335
rect 10 3310 40 3315
rect 10 3235 40 3240
rect 10 3215 15 3235
rect 15 3215 35 3235
rect 35 3215 40 3235
rect 10 3210 40 3215
rect 10 3135 40 3140
rect 10 3115 15 3135
rect 15 3115 35 3135
rect 35 3115 40 3135
rect 10 3110 40 3115
rect 210 3535 240 3540
rect 210 3515 215 3535
rect 215 3515 235 3535
rect 235 3515 240 3535
rect 210 3510 240 3515
rect 210 3435 240 3440
rect 210 3415 215 3435
rect 215 3415 235 3435
rect 235 3415 240 3435
rect 210 3410 240 3415
rect 210 3335 240 3340
rect 210 3315 215 3335
rect 215 3315 235 3335
rect 235 3315 240 3335
rect 210 3310 240 3315
rect 210 3235 240 3240
rect 210 3215 215 3235
rect 215 3215 235 3235
rect 235 3215 240 3235
rect 210 3210 240 3215
rect 110 3035 140 3040
rect 110 3015 115 3035
rect 115 3015 135 3035
rect 135 3015 140 3035
rect 110 3010 140 3015
rect 10 2810 40 2840
rect 210 2810 240 2840
rect 10 2435 40 2440
rect 10 2415 15 2435
rect 15 2415 35 2435
rect 35 2415 40 2435
rect 10 2410 40 2415
rect 10 2335 40 2340
rect 10 2315 15 2335
rect 15 2315 35 2335
rect 35 2315 40 2335
rect 10 2310 40 2315
rect 10 2235 40 2240
rect 10 2215 15 2235
rect 15 2215 35 2235
rect 35 2215 40 2235
rect 10 2210 40 2215
rect 10 2135 40 2140
rect 10 2115 15 2135
rect 15 2115 35 2135
rect 35 2115 40 2135
rect 10 2110 40 2115
rect 10 2035 40 2040
rect 10 2015 15 2035
rect 15 2015 35 2035
rect 35 2015 40 2035
rect 10 2010 40 2015
rect 10 1835 40 1840
rect 10 1815 15 1835
rect 15 1815 35 1835
rect 35 1815 40 1835
rect 10 1810 40 1815
rect 10 1735 40 1740
rect 10 1715 15 1735
rect 15 1715 35 1735
rect 35 1715 40 1735
rect 10 1710 40 1715
rect 10 1635 40 1640
rect 10 1615 15 1635
rect 15 1615 35 1635
rect 35 1615 40 1635
rect 10 1610 40 1615
rect 10 1535 40 1540
rect 10 1515 15 1535
rect 15 1515 35 1535
rect 35 1515 40 1535
rect 10 1510 40 1515
rect 10 1435 40 1440
rect 10 1415 15 1435
rect 15 1415 35 1435
rect 35 1415 40 1435
rect 10 1410 40 1415
rect 110 1935 140 1940
rect 110 1915 115 1935
rect 115 1915 135 1935
rect 135 1915 140 1935
rect 110 1910 140 1915
rect 210 2435 240 2440
rect 210 2415 215 2435
rect 215 2415 235 2435
rect 235 2415 240 2435
rect 210 2410 240 2415
rect 210 2335 240 2340
rect 210 2315 215 2335
rect 215 2315 235 2335
rect 235 2315 240 2335
rect 210 2310 240 2315
rect 210 2235 240 2240
rect 210 2215 215 2235
rect 215 2215 235 2235
rect 235 2215 240 2235
rect 210 2210 240 2215
rect 210 2135 240 2140
rect 210 2115 215 2135
rect 215 2115 235 2135
rect 235 2115 240 2135
rect 210 2110 240 2115
rect 210 2035 240 2040
rect 210 2015 215 2035
rect 215 2015 235 2035
rect 235 2015 240 2035
rect 210 2010 240 2015
rect 210 1835 240 1840
rect 210 1815 215 1835
rect 215 1815 235 1835
rect 235 1815 240 1835
rect 210 1810 240 1815
rect 210 1735 240 1740
rect 210 1715 215 1735
rect 215 1715 235 1735
rect 235 1715 240 1735
rect 210 1710 240 1715
rect 210 1635 240 1640
rect 210 1615 215 1635
rect 215 1615 235 1635
rect 235 1615 240 1635
rect 210 1610 240 1615
rect 210 1535 240 1540
rect 210 1515 215 1535
rect 215 1515 235 1535
rect 235 1515 240 1535
rect 210 1510 240 1515
rect 210 1435 240 1440
rect 210 1415 215 1435
rect 215 1415 235 1435
rect 235 1415 240 1435
rect 210 1410 240 1415
rect 10 1010 40 1040
rect 210 1010 240 1040
rect 110 835 140 840
rect 110 815 115 835
rect 115 815 135 835
rect 135 815 140 835
rect 110 810 140 815
rect 10 735 40 740
rect 10 715 15 735
rect 15 715 35 735
rect 35 715 40 735
rect 10 710 40 715
rect 10 635 40 640
rect 10 615 15 635
rect 15 615 35 635
rect 35 615 40 635
rect 10 610 40 615
rect 10 535 40 540
rect 10 515 15 535
rect 15 515 35 535
rect 35 515 40 535
rect 10 510 40 515
rect 10 435 40 440
rect 10 415 15 435
rect 15 415 35 435
rect 35 415 40 435
rect 10 410 40 415
rect 10 335 40 340
rect 10 315 15 335
rect 15 315 35 335
rect 35 315 40 335
rect 10 310 40 315
rect 210 635 240 640
rect 210 615 215 635
rect 215 615 235 635
rect 235 615 240 635
rect 210 610 240 615
rect 210 535 240 540
rect 210 515 215 535
rect 215 515 235 535
rect 235 515 240 535
rect 210 510 240 515
rect 210 435 240 440
rect 210 415 215 435
rect 215 415 235 435
rect 235 415 240 435
rect 210 410 240 415
rect 210 335 240 340
rect 210 315 215 335
rect 215 315 235 335
rect 235 315 240 335
rect 210 310 240 315
rect 10 210 40 240
rect 10 110 40 140
rect 210 210 240 240
rect 210 110 240 140
<< metal2 >>
rect 0 3740 250 3750
rect 0 3710 10 3740
rect 40 3710 210 3740
rect 240 3710 250 3740
rect 0 3700 250 3710
rect 0 3640 250 3650
rect 0 3610 10 3640
rect 40 3610 210 3640
rect 240 3610 250 3640
rect 0 3600 250 3610
rect 0 3540 250 3550
rect 0 3510 10 3540
rect 40 3510 210 3540
rect 240 3510 250 3540
rect 0 3500 250 3510
rect 0 3440 250 3450
rect 0 3410 10 3440
rect 40 3410 210 3440
rect 240 3410 250 3440
rect 0 3400 250 3410
rect 0 3340 250 3350
rect 0 3310 10 3340
rect 40 3310 210 3340
rect 240 3310 250 3340
rect 0 3300 250 3310
rect 0 3240 250 3250
rect 0 3210 10 3240
rect 40 3210 210 3240
rect 240 3210 250 3240
rect 0 3200 250 3210
rect 0 3140 250 3150
rect 0 3110 10 3140
rect 40 3110 210 3140
rect 240 3110 250 3140
rect 0 3100 250 3110
rect 100 3040 150 3050
rect 100 3010 110 3040
rect 140 3010 150 3040
rect 100 3000 150 3010
rect 0 2840 250 2850
rect 0 2810 10 2840
rect 40 2810 210 2840
rect 240 2810 250 2840
rect 0 2800 250 2810
rect 0 2440 250 2450
rect 0 2410 10 2440
rect 40 2410 210 2440
rect 240 2410 250 2440
rect 0 2400 250 2410
rect 0 2340 250 2350
rect 0 2310 10 2340
rect 40 2310 210 2340
rect 240 2310 250 2340
rect 0 2300 250 2310
rect 0 2240 250 2250
rect 0 2210 10 2240
rect 40 2210 210 2240
rect 240 2210 250 2240
rect 0 2200 250 2210
rect 0 2140 250 2150
rect 0 2110 10 2140
rect 40 2110 210 2140
rect 240 2110 250 2140
rect 0 2100 250 2110
rect 0 2040 250 2050
rect 0 2010 10 2040
rect 40 2010 210 2040
rect 240 2010 250 2040
rect 0 2000 250 2010
rect 100 1940 150 1950
rect 100 1910 110 1940
rect 140 1910 150 1940
rect 100 1900 150 1910
rect 0 1840 250 1850
rect 0 1810 10 1840
rect 40 1810 210 1840
rect 240 1810 250 1840
rect 0 1800 250 1810
rect 0 1740 250 1750
rect 0 1710 10 1740
rect 40 1710 210 1740
rect 240 1710 250 1740
rect 0 1700 250 1710
rect 0 1640 250 1650
rect 0 1610 10 1640
rect 40 1610 210 1640
rect 240 1610 250 1640
rect 0 1600 250 1610
rect 0 1540 250 1550
rect 0 1510 10 1540
rect 40 1510 210 1540
rect 240 1510 250 1540
rect 0 1500 250 1510
rect 0 1440 250 1450
rect 0 1410 10 1440
rect 40 1410 210 1440
rect 240 1410 250 1440
rect 0 1400 250 1410
rect 0 1040 250 1050
rect 0 1010 10 1040
rect 40 1010 210 1040
rect 240 1010 250 1040
rect 0 1000 250 1010
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 100 800 150 810
rect 0 740 250 750
rect 0 710 10 740
rect 40 710 210 740
rect 240 710 250 740
rect 0 700 250 710
rect 0 640 250 650
rect 0 610 10 640
rect 40 610 210 640
rect 240 610 250 640
rect 0 600 250 610
rect 0 540 250 550
rect 0 510 10 540
rect 40 510 210 540
rect 240 510 250 540
rect 0 500 250 510
rect 0 440 250 450
rect 0 410 10 440
rect 40 410 210 440
rect 240 410 250 440
rect 0 400 250 410
rect 0 340 250 350
rect 0 310 10 340
rect 40 310 210 340
rect 240 310 250 340
rect 0 300 250 310
rect 0 240 250 250
rect 0 210 10 240
rect 40 210 210 240
rect 240 210 250 240
rect 0 200 250 210
rect 0 140 250 150
rect 0 110 10 140
rect 40 110 210 140
rect 240 110 250 140
rect 0 100 250 110
<< via2 >>
rect 10 3710 40 3740
rect 210 3710 240 3740
rect 10 3610 40 3640
rect 210 3610 240 3640
rect 10 3510 40 3540
rect 210 3510 240 3540
rect 10 3410 40 3440
rect 210 3410 240 3440
rect 10 3310 40 3340
rect 210 3310 240 3340
rect 10 3210 40 3240
rect 210 3210 240 3240
rect 10 3110 40 3140
rect 210 3110 240 3140
rect 110 3010 140 3040
rect 10 2810 40 2840
rect 210 2810 240 2840
rect 10 2410 40 2440
rect 210 2410 240 2440
rect 10 2210 40 2240
rect 210 2210 240 2240
rect 10 2010 40 2040
rect 210 2010 240 2040
rect 110 1910 140 1940
rect 10 1810 40 1840
rect 210 1810 240 1840
rect 10 1610 40 1640
rect 210 1610 240 1640
rect 10 1410 40 1440
rect 210 1410 240 1440
rect 10 1010 40 1040
rect 210 1010 240 1040
rect 110 810 140 840
rect 10 710 40 740
rect 210 710 240 740
rect 10 610 40 640
rect 210 610 240 640
rect 10 510 40 540
rect 210 510 240 540
rect 10 410 40 440
rect 210 410 240 440
rect 10 310 40 340
rect 210 310 240 340
rect 10 210 40 240
rect 210 210 240 240
rect 10 110 40 140
rect 210 110 240 140
<< metal3 >>
rect 0 3740 250 3750
rect 0 3710 10 3740
rect 40 3710 210 3740
rect 240 3710 250 3740
rect 0 3700 250 3710
rect 0 3640 250 3650
rect 0 3610 10 3640
rect 40 3610 210 3640
rect 240 3610 250 3640
rect 0 3600 250 3610
rect 0 3540 250 3550
rect 0 3510 10 3540
rect 40 3510 210 3540
rect 240 3510 250 3540
rect 0 3500 250 3510
rect 0 3440 250 3450
rect 0 3410 10 3440
rect 40 3410 210 3440
rect 240 3410 250 3440
rect 0 3400 250 3410
rect 0 3340 250 3350
rect 0 3310 10 3340
rect 40 3310 210 3340
rect 240 3310 250 3340
rect 0 3300 250 3310
rect 0 3240 250 3250
rect 0 3210 10 3240
rect 40 3210 210 3240
rect 240 3210 250 3240
rect 0 3200 250 3210
rect 0 3140 250 3150
rect 0 3110 10 3140
rect 40 3110 210 3140
rect 240 3110 250 3140
rect 0 3100 250 3110
rect 100 3040 150 3050
rect 100 3010 110 3040
rect 140 3010 150 3040
rect 100 3000 150 3010
rect 0 2840 250 2850
rect 0 2810 10 2840
rect 40 2810 210 2840
rect 240 2810 250 2840
rect 0 2800 250 2810
rect 0 2440 250 2450
rect 0 2410 10 2440
rect 40 2410 210 2440
rect 240 2410 250 2440
rect 0 2400 250 2410
rect 0 2240 250 2250
rect 0 2210 10 2240
rect 40 2210 210 2240
rect 240 2210 250 2240
rect 0 2200 250 2210
rect 0 2040 250 2050
rect 0 2010 10 2040
rect 40 2010 210 2040
rect 240 2010 250 2040
rect 0 2000 250 2010
rect 100 1940 150 1950
rect 100 1910 110 1940
rect 140 1910 150 1940
rect 100 1900 150 1910
rect 0 1840 250 1850
rect 0 1810 10 1840
rect 40 1810 210 1840
rect 240 1810 250 1840
rect 0 1800 250 1810
rect 0 1640 250 1650
rect 0 1610 10 1640
rect 40 1610 210 1640
rect 240 1610 250 1640
rect 0 1600 250 1610
rect 0 1440 250 1450
rect 0 1410 10 1440
rect 40 1410 210 1440
rect 240 1410 250 1440
rect 0 1400 250 1410
rect 0 1040 250 1050
rect 0 1010 10 1040
rect 40 1010 210 1040
rect 240 1010 250 1040
rect 0 1000 250 1010
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 100 800 150 810
rect 0 740 250 750
rect 0 710 10 740
rect 40 710 210 740
rect 240 710 250 740
rect 0 700 250 710
rect 0 640 250 650
rect 0 610 10 640
rect 40 610 210 640
rect 240 610 250 640
rect 0 600 250 610
rect 0 540 250 550
rect 0 510 10 540
rect 40 510 210 540
rect 240 510 250 540
rect 0 500 250 510
rect 0 440 250 450
rect 0 410 10 440
rect 40 410 210 440
rect 240 410 250 440
rect 0 400 250 410
rect 0 340 250 350
rect 0 310 10 340
rect 40 310 210 340
rect 240 310 250 340
rect 0 300 250 310
rect 0 240 250 250
rect 0 210 10 240
rect 40 210 210 240
rect 240 210 250 240
rect 0 200 250 210
rect 0 140 250 150
rect 0 110 10 140
rect 40 110 210 140
rect 240 110 250 140
rect 0 100 250 110
<< labels >>
rlabel locali 0 2900 250 2950 0 bp
port 3 nsew
rlabel locali 0 900 250 950 0 bp
port 3 nsew
rlabel locali 50 2750 200 2800 0 bn
port 4 nsew
rlabel locali 50 1050 200 1100 0 bn
port 4 nsew
rlabel metal3 50 3700 200 3750 0 vdd
port 5 nsew
rlabel metal3 50 2800 200 2850 0 vss
port 6 nsew
rlabel metal3 50 1000 200 1050 0 vss
port 6 nsew
rlabel locali 0 3800 300 3850 0 vsub
port 7 nsew
rlabel locali 0 0 300 50 0 vsub
port 7 nsew
rlabel metal3 50 100 200 150 0 vdd
port 5 nsew
rlabel metal1 100 1950 150 2000 0 xn
rlabel metal1 100 3050 150 3100 0 xpt
rlabel metal1 100 750 150 800 0 xpb
<< end >>
