magic
tech sky130A
timestamp 1726841226
<< pwell >>
rect 2300 2500 2350 2750
rect 4550 2500 4600 2750
rect 5900 2500 5950 2750
rect 6350 2500 6400 2750
rect 500 2100 550 2150
rect 3200 2100 3250 2150
rect 4100 1700 4150 1750
rect 6800 1700 6850 1750
rect 950 1200 1000 1350
rect 1400 1200 1450 1350
rect 2750 1100 2800 1350
rect 5000 1100 5050 1350
<< locali >>
rect 50 3800 7300 3850
rect 50 2900 7300 2950
rect 50 2750 7300 2800
rect 50 1050 7300 1100
rect 50 900 7300 950
rect 50 0 7300 50
<< metal1 >>
rect 4550 2740 4600 2750
rect 4550 2710 4560 2740
rect 4590 2710 4600 2740
rect 4550 2690 4600 2710
rect 4550 2660 4560 2690
rect 4590 2660 4600 2690
rect 4550 2640 4600 2660
rect 4550 2610 4560 2640
rect 4590 2610 4600 2640
rect 4550 2590 4600 2610
rect 4550 2560 4560 2590
rect 4590 2560 4600 2590
rect 4550 2540 4600 2560
rect 4550 2510 4560 2540
rect 4590 2510 4600 2540
rect 4550 2500 4600 2510
rect 6350 2740 6400 2750
rect 6350 2710 6360 2740
rect 6390 2710 6400 2740
rect 6350 2690 6400 2710
rect 6350 2660 6360 2690
rect 6390 2660 6400 2690
rect 6350 2640 6400 2660
rect 6350 2610 6360 2640
rect 6390 2610 6400 2640
rect 6350 2590 6400 2610
rect 6350 2560 6360 2590
rect 6390 2560 6400 2590
rect 6350 2540 6400 2560
rect 6350 2510 6360 2540
rect 6390 2510 6400 2540
rect 6350 2500 6400 2510
rect 950 1340 1000 1350
rect 950 1310 960 1340
rect 990 1310 1000 1340
rect 950 1290 1000 1310
rect 950 1260 960 1290
rect 990 1260 1000 1290
rect 950 1240 1000 1260
rect 950 1210 960 1240
rect 990 1210 1000 1240
rect 950 1190 1000 1210
rect 950 1160 960 1190
rect 990 1160 1000 1190
rect 950 1140 1000 1160
rect 950 1110 960 1140
rect 990 1110 1000 1140
rect 950 1100 1000 1110
rect 2750 1340 2800 1350
rect 2750 1310 2760 1340
rect 2790 1310 2800 1340
rect 2750 1290 2800 1310
rect 2750 1260 2760 1290
rect 2790 1260 2800 1290
rect 2750 1240 2800 1260
rect 2750 1210 2760 1240
rect 2790 1210 2800 1240
rect 2750 1190 2800 1210
rect 2750 1160 2760 1190
rect 2790 1160 2800 1190
rect 2750 1140 2800 1160
rect 2750 1110 2760 1140
rect 2790 1110 2800 1140
rect 2750 1100 2800 1110
<< via1 >>
rect 4560 2710 4590 2740
rect 4560 2660 4590 2690
rect 4560 2610 4590 2640
rect 4560 2560 4590 2590
rect 4560 2510 4590 2540
rect 6360 2710 6390 2740
rect 6360 2660 6390 2690
rect 6360 2610 6390 2640
rect 6360 2560 6390 2590
rect 6360 2510 6390 2540
rect 960 1310 990 1340
rect 960 1260 990 1290
rect 960 1210 990 1240
rect 960 1160 990 1190
rect 960 1110 990 1140
rect 2760 1310 2790 1340
rect 2760 1260 2790 1290
rect 2760 1210 2790 1240
rect 2760 1160 2790 1190
rect 2760 1110 2790 1140
<< metal2 >>
rect 4550 2740 4600 2750
rect 4550 2710 4560 2740
rect 4590 2710 4600 2740
rect 4550 2690 4600 2710
rect 4550 2660 4560 2690
rect 4590 2660 4600 2690
rect 4550 2640 4600 2660
rect 4550 2610 4560 2640
rect 4590 2610 4600 2640
rect 4550 2590 4600 2610
rect 4550 2560 4560 2590
rect 4590 2560 4600 2590
rect 4550 2540 4600 2560
rect 4550 2510 4560 2540
rect 4590 2510 4600 2540
rect 4550 2500 4600 2510
rect 6350 2740 6400 2750
rect 6350 2710 6360 2740
rect 6390 2710 6400 2740
rect 6350 2690 6400 2710
rect 6350 2660 6360 2690
rect 6390 2660 6400 2690
rect 6350 2640 6400 2660
rect 6350 2610 6360 2640
rect 6390 2610 6400 2640
rect 6350 2590 6400 2610
rect 6350 2560 6360 2590
rect 6390 2560 6400 2590
rect 6350 2540 6400 2560
rect 6350 2510 6360 2540
rect 6390 2510 6400 2540
rect 6350 2500 6400 2510
rect 950 1340 1000 1350
rect 950 1310 960 1340
rect 990 1310 1000 1340
rect 950 1290 1000 1310
rect 950 1260 960 1290
rect 990 1260 1000 1290
rect 950 1240 1000 1260
rect 950 1210 960 1240
rect 990 1210 1000 1240
rect 950 1190 1000 1210
rect 950 1160 960 1190
rect 990 1160 1000 1190
rect 950 1140 1000 1160
rect 950 1110 960 1140
rect 990 1110 1000 1140
rect 950 1100 1000 1110
rect 2750 1340 2800 1350
rect 2750 1310 2760 1340
rect 2790 1310 2800 1340
rect 2750 1290 2800 1310
rect 2750 1260 2760 1290
rect 2790 1260 2800 1290
rect 2750 1240 2800 1260
rect 2750 1210 2760 1240
rect 2790 1210 2800 1240
rect 2750 1190 2800 1210
rect 2750 1160 2760 1190
rect 2790 1160 2800 1190
rect 2750 1140 2800 1160
rect 2750 1110 2760 1140
rect 2790 1110 2800 1140
rect 2750 1100 2800 1110
<< via2 >>
rect 4560 2710 4590 2740
rect 4560 2660 4590 2690
rect 4560 2610 4590 2640
rect 4560 2560 4590 2590
rect 4560 2510 4590 2540
rect 6360 2710 6390 2740
rect 6360 2660 6390 2690
rect 6360 2610 6390 2640
rect 6360 2560 6390 2590
rect 6360 2510 6390 2540
rect 960 1310 990 1340
rect 960 1260 990 1290
rect 960 1210 990 1240
rect 960 1160 990 1190
rect 960 1110 990 1140
rect 2760 1310 2790 1340
rect 2760 1260 2790 1290
rect 2760 1210 2790 1240
rect 2760 1160 2790 1190
rect 2760 1110 2790 1140
<< metal3 >>
rect 50 3700 7300 3750
rect 50 2800 7300 2850
rect 50 2745 7300 2750
rect 50 2705 2305 2745
rect 2345 2740 5905 2745
rect 2345 2710 4560 2740
rect 4590 2710 5905 2740
rect 2345 2705 5905 2710
rect 5945 2740 7300 2745
rect 5945 2710 6360 2740
rect 6390 2710 7300 2740
rect 5945 2705 7300 2710
rect 50 2695 7300 2705
rect 50 2655 2305 2695
rect 2345 2690 5905 2695
rect 2345 2660 4560 2690
rect 4590 2660 5905 2690
rect 2345 2655 5905 2660
rect 5945 2690 7300 2695
rect 5945 2660 6360 2690
rect 6390 2660 7300 2690
rect 5945 2655 7300 2660
rect 50 2645 7300 2655
rect 50 2605 2305 2645
rect 2345 2640 5905 2645
rect 2345 2610 4560 2640
rect 4590 2610 5905 2640
rect 2345 2605 5905 2610
rect 5945 2640 7300 2645
rect 5945 2610 6360 2640
rect 6390 2610 7300 2640
rect 5945 2605 7300 2610
rect 50 2595 7300 2605
rect 50 2555 2305 2595
rect 2345 2590 5905 2595
rect 2345 2560 4560 2590
rect 4590 2560 5905 2590
rect 2345 2555 5905 2560
rect 5945 2590 7300 2595
rect 5945 2560 6360 2590
rect 6390 2560 7300 2590
rect 5945 2555 7300 2560
rect 50 2545 7300 2555
rect 50 2505 2305 2545
rect 2345 2540 5905 2545
rect 2345 2510 4560 2540
rect 4590 2510 5905 2540
rect 2345 2505 5905 2510
rect 5945 2540 7300 2545
rect 5945 2510 6360 2540
rect 6390 2510 7300 2540
rect 5945 2505 7300 2510
rect 50 2500 7300 2505
rect 50 2145 7300 2150
rect 50 2105 505 2145
rect 545 2105 3205 2145
rect 3245 2105 7300 2145
rect 50 2100 7300 2105
rect 50 1745 7300 1750
rect 50 1705 4105 1745
rect 4145 1705 6805 1745
rect 6845 1705 7300 1745
rect 50 1700 7300 1705
rect 50 1345 7300 1350
rect 50 1340 1405 1345
rect 50 1310 960 1340
rect 990 1310 1405 1340
rect 50 1305 1405 1310
rect 1445 1340 5005 1345
rect 1445 1310 2760 1340
rect 2790 1310 5005 1340
rect 1445 1305 5005 1310
rect 5045 1305 7300 1345
rect 50 1295 7300 1305
rect 50 1290 1405 1295
rect 50 1260 960 1290
rect 990 1260 1405 1290
rect 50 1255 1405 1260
rect 1445 1290 5005 1295
rect 1445 1260 2760 1290
rect 2790 1260 5005 1290
rect 1445 1255 5005 1260
rect 5045 1255 7300 1295
rect 50 1245 7300 1255
rect 50 1240 1405 1245
rect 50 1210 960 1240
rect 990 1210 1405 1240
rect 50 1205 1405 1210
rect 1445 1240 5005 1245
rect 1445 1210 2760 1240
rect 2790 1210 5005 1240
rect 1445 1205 5005 1210
rect 5045 1205 7300 1245
rect 50 1195 7300 1205
rect 50 1190 1405 1195
rect 50 1160 960 1190
rect 990 1160 1405 1190
rect 50 1155 1405 1160
rect 1445 1190 5005 1195
rect 1445 1160 2760 1190
rect 2790 1160 5005 1190
rect 1445 1155 5005 1160
rect 5045 1155 7300 1195
rect 50 1145 7300 1155
rect 50 1140 1405 1145
rect 50 1110 960 1140
rect 990 1110 1405 1140
rect 50 1105 1405 1110
rect 1445 1140 5005 1145
rect 1445 1110 2760 1140
rect 2790 1110 5005 1140
rect 1445 1105 5005 1110
rect 5045 1105 7300 1145
rect 50 1100 7300 1105
rect 50 1000 7300 1050
rect 50 100 7300 150
<< via3 >>
rect 2305 2705 2345 2745
rect 5905 2705 5945 2745
rect 2305 2655 2345 2695
rect 5905 2655 5945 2695
rect 2305 2605 2345 2645
rect 5905 2605 5945 2645
rect 2305 2555 2345 2595
rect 5905 2555 5945 2595
rect 2305 2505 2345 2545
rect 5905 2505 5945 2545
rect 505 2105 545 2145
rect 3205 2105 3245 2145
rect 4105 1705 4145 1745
rect 6805 1705 6845 1745
rect 1405 1305 1445 1345
rect 5005 1305 5045 1345
rect 1405 1255 1445 1295
rect 5005 1255 5045 1295
rect 1405 1205 1445 1245
rect 5005 1205 5045 1245
rect 1405 1155 1445 1195
rect 5005 1155 5045 1195
rect 1405 1105 1445 1145
rect 5005 1105 5045 1145
<< metal4 >>
rect 2300 2745 2350 2750
rect 2300 2705 2305 2745
rect 2345 2705 2350 2745
rect 2300 2695 2350 2705
rect 2300 2655 2305 2695
rect 2345 2655 2350 2695
rect 2300 2645 2350 2655
rect 2300 2605 2305 2645
rect 2345 2605 2350 2645
rect 2300 2595 2350 2605
rect 2300 2555 2305 2595
rect 2345 2555 2350 2595
rect 2300 2545 2350 2555
rect 2300 2505 2305 2545
rect 2345 2505 2350 2545
rect 2300 2500 2350 2505
rect 5900 2745 5950 2750
rect 5900 2705 5905 2745
rect 5945 2705 5950 2745
rect 5900 2695 5950 2705
rect 5900 2655 5905 2695
rect 5945 2655 5950 2695
rect 5900 2645 5950 2655
rect 5900 2605 5905 2645
rect 5945 2605 5950 2645
rect 5900 2595 5950 2605
rect 5900 2555 5905 2595
rect 5945 2555 5950 2595
rect 5900 2545 5950 2555
rect 5900 2505 5905 2545
rect 5945 2505 5950 2545
rect 5900 2500 5950 2505
rect 500 2145 550 2150
rect 500 2105 505 2145
rect 545 2105 550 2145
rect 500 2100 550 2105
rect 3200 2145 3250 2150
rect 3200 2105 3205 2145
rect 3245 2105 3250 2145
rect 3200 2100 3250 2105
rect 4100 1745 4150 1750
rect 4100 1705 4105 1745
rect 4145 1705 4150 1745
rect 4100 1700 4150 1705
rect 6800 1745 6850 1750
rect 6800 1705 6805 1745
rect 6845 1705 6850 1745
rect 6800 1700 6850 1705
rect 1400 1345 1450 1350
rect 1400 1305 1405 1345
rect 1445 1305 1450 1345
rect 1400 1295 1450 1305
rect 1400 1255 1405 1295
rect 1445 1255 1450 1295
rect 1400 1245 1450 1255
rect 1400 1205 1405 1245
rect 1445 1205 1450 1245
rect 1400 1195 1450 1205
rect 1400 1155 1405 1195
rect 1445 1155 1450 1195
rect 1400 1145 1450 1155
rect 1400 1105 1405 1145
rect 1445 1105 1450 1145
rect 1400 1100 1450 1105
rect 5000 1345 5050 1350
rect 5000 1305 5005 1345
rect 5045 1305 5050 1345
rect 5000 1295 5050 1305
rect 5000 1255 5005 1295
rect 5045 1255 5050 1295
rect 5000 1245 5050 1255
rect 5000 1205 5005 1245
rect 5045 1205 5050 1245
rect 5000 1195 5050 1205
rect 5000 1155 5005 1195
rect 5045 1155 5050 1195
rect 5000 1145 5050 1155
rect 5000 1105 5005 1145
rect 5045 1105 5050 1145
rect 5000 1100 5050 1105
use inv1p1  a0
timestamp 1726000395
transform 1 0 50 0 1 0
box -50 0 1000 3850
use inv1p1  a1
timestamp 1726000395
transform -1 0 1900 0 1 0
box -50 0 1000 3850
use inv1p1  a2
timestamp 1726000395
transform 1 0 1850 0 1 0
box -50 0 1000 3850
use inv1p1  a3
timestamp 1726000395
transform -1 0 3700 0 1 0
box -50 0 1000 3850
use inv1p1  a4
timestamp 1726000395
transform 1 0 3650 0 1 0
box -50 0 1000 3850
use inv1p1  a5
timestamp 1726000395
transform -1 0 5500 0 1 0
box -50 0 1000 3850
use inv1p1  a6
timestamp 1726000395
transform 1 0 5450 0 1 0
box -50 0 1000 3850
use inv1p1  a7
timestamp 1726000395
transform -1 0 7300 0 1 0
box -50 0 1000 3850
<< labels >>
rlabel metal3 50 2100 7300 2150 0 ip
port 1 nsew
rlabel metal3 50 1700 7300 1750 0 im
port 2 nsew
rlabel metal3 50 2500 7300 2750 0 op
port 5 nsew
rlabel metal3 50 1100 7300 1350 0 om
port 6 nsew
rlabel locali 50 2900 7300 2950 0 bp
port 7 nsew
rlabel locali 50 900 7300 950 0 bp
port 7 nsew
rlabel locali 50 2750 7300 2800 0 bn
port 8 nsew
rlabel locali 50 1050 7300 1100 0 bn
port 8 nsew
rlabel metal3 50 3700 7300 3750 0 vreg
port 9 nsew
rlabel metal3 50 100 7300 150 0 vreg
port 9 nsew
rlabel metal3 50 2800 7300 2850 0 vss
port 10 nsew
rlabel metal3 50 1000 7300 1050 0 vss
port 10 nsew
rlabel locali 50 3800 7300 3850 0 vsub
port 11 nsew
rlabel locali 50 0 7300 50 0 vsub
port 11 nsew
<< end >>
