magic
tech sky130A
timestamp 1719349916
<< error_s >>
rect 2700 2300 3150 2750
rect -200 900 250 1350
<< dnwell >>
rect -200 750 3150 2900
<< nwell >>
rect -200 3550 -150 3600
<< mvndiffc >>
rect 2465 2515 2485 2535
rect 2865 2515 2885 2535
<< locali >>
rect -200 3700 3150 3750
rect -200 3550 3050 3600
rect -200 50 3050 100
rect -200 -100 3150 -50
<< viali >>
rect 865 2515 885 2535
rect 1265 2515 1285 2535
rect 2465 2515 2485 2535
rect 2865 2515 2885 2535
rect 465 1115 485 1135
rect 1665 1115 1685 1135
rect 2065 1115 2085 1135
<< metal1 >>
rect 850 2540 900 2550
rect 850 2510 860 2540
rect 890 2510 900 2540
rect 850 2500 900 2510
rect 1250 2540 1300 2550
rect 1250 2510 1260 2540
rect 1290 2510 1300 2540
rect 1250 2500 1300 2510
rect 2450 2540 2500 2550
rect 2450 2510 2460 2540
rect 2490 2510 2500 2540
rect 2450 2500 2500 2510
rect 2850 2540 2900 2550
rect 2850 2510 2860 2540
rect 2890 2510 2900 2540
rect 2850 2500 2900 2510
rect 450 1140 500 1150
rect 450 1110 460 1140
rect 490 1110 500 1140
rect 450 1100 500 1110
rect 1650 1140 1700 1150
rect 1650 1110 1660 1140
rect 1690 1110 1700 1140
rect 1650 1100 1700 1110
rect 2050 1140 2100 1150
rect 2050 1110 2060 1140
rect 2090 1110 2100 1140
rect 2050 1100 2100 1110
<< via1 >>
rect 860 2535 890 2540
rect 860 2515 865 2535
rect 865 2515 885 2535
rect 885 2515 890 2535
rect 860 2510 890 2515
rect 1260 2535 1290 2540
rect 1260 2515 1265 2535
rect 1265 2515 1285 2535
rect 1285 2515 1290 2535
rect 1260 2510 1290 2515
rect 2460 2535 2490 2540
rect 2460 2515 2465 2535
rect 2465 2515 2485 2535
rect 2485 2515 2490 2535
rect 2460 2510 2490 2515
rect 2860 2535 2890 2540
rect 2860 2515 2865 2535
rect 2865 2515 2885 2535
rect 2885 2515 2890 2535
rect 2860 2510 2890 2515
rect 60 1110 90 1140
rect 460 1135 490 1140
rect 460 1115 465 1135
rect 465 1115 485 1135
rect 485 1115 490 1135
rect 460 1110 490 1115
rect 1660 1135 1690 1140
rect 1660 1115 1665 1135
rect 1665 1115 1685 1135
rect 1685 1115 1690 1135
rect 1660 1110 1690 1115
rect 2060 1135 2090 1140
rect 2060 1115 2065 1135
rect 2065 1115 2085 1135
rect 2085 1115 2090 1135
rect 2060 1110 2090 1115
<< metal2 >>
rect 850 2540 900 2550
rect 850 2510 860 2540
rect 890 2510 900 2540
rect 850 2500 900 2510
rect 1250 2540 1300 2550
rect 1250 2510 1260 2540
rect 1290 2510 1300 2540
rect 1250 2500 1300 2510
rect 2450 2540 2500 2550
rect 2450 2510 2460 2540
rect 2490 2510 2500 2540
rect 2450 2500 2500 2510
rect 2850 2540 2900 2550
rect 2850 2510 2860 2540
rect 2890 2510 2900 2540
rect 2850 2500 2900 2510
rect 2350 2200 2400 2250
rect 2950 2200 3000 2250
rect 1550 2000 1600 2050
rect 2150 2000 2200 2050
rect 50 1140 100 1150
rect 50 1110 60 1140
rect 90 1110 100 1140
rect 50 1100 100 1110
rect 450 1140 500 1150
rect 450 1110 460 1140
rect 490 1110 500 1140
rect 450 1100 500 1110
rect 1650 1140 1700 1150
rect 1650 1110 1660 1140
rect 1690 1110 1700 1140
rect 1650 1100 1700 1110
rect 2050 1140 2100 1150
rect 2050 1110 2060 1140
rect 2090 1110 2100 1140
rect 2050 1100 2100 1110
<< via2 >>
rect 860 2510 890 2540
rect 1260 2510 1290 2540
rect 2460 2510 2490 2540
rect 2860 2510 2890 2540
rect 60 1110 90 1140
rect 460 1110 490 1140
rect 1660 1110 1690 1140
rect 2060 1110 2090 1140
<< metal3 >>
rect -200 3400 -100 3450
rect -150 2700 3100 2750
rect -150 2545 3100 2650
rect -150 2505 355 2545
rect 395 2540 955 2545
rect 395 2510 860 2540
rect 890 2510 955 2540
rect 395 2505 955 2510
rect 995 2540 1955 2545
rect 995 2510 1260 2540
rect 1290 2510 1955 2540
rect 995 2505 1955 2510
rect 1995 2540 2555 2545
rect 1995 2510 2460 2540
rect 2490 2510 2555 2540
rect 1995 2505 2555 2510
rect 2595 2540 3100 2545
rect 2595 2510 2860 2540
rect 2890 2510 3100 2540
rect 2595 2505 3100 2510
rect -150 2400 3100 2505
rect -150 2245 3100 2250
rect -150 2205 2355 2245
rect 2395 2205 2955 2245
rect 2995 2205 3100 2245
rect -150 2200 3100 2205
rect -150 2045 3100 2050
rect -150 2005 1555 2045
rect 1595 2005 2155 2045
rect 2195 2005 3100 2045
rect -150 2000 3100 2005
rect -150 1645 3100 1650
rect -150 1605 -45 1645
rect -5 1605 555 1645
rect 595 1605 3100 1645
rect -150 1600 3100 1605
rect -150 1445 3100 1450
rect -150 1405 755 1445
rect 795 1405 1355 1445
rect 1395 1405 3100 1445
rect -150 1400 3100 1405
rect -150 1145 3100 1250
rect -150 1140 155 1145
rect -150 1110 60 1140
rect 90 1110 155 1140
rect -150 1105 155 1110
rect 195 1140 1155 1145
rect 195 1110 460 1140
rect 490 1110 1155 1140
rect 195 1105 1155 1110
rect 1195 1140 1755 1145
rect 1195 1110 1660 1140
rect 1690 1110 1755 1140
rect 1195 1105 1755 1110
rect 1795 1140 2755 1145
rect 1795 1110 2060 1140
rect 2090 1110 2755 1140
rect 1795 1105 2755 1110
rect 2795 1105 3100 1145
rect -150 1000 3100 1105
rect -150 900 3100 950
rect -200 200 -150 250
<< via3 >>
rect 355 2505 395 2545
rect 955 2505 995 2545
rect 1955 2505 1995 2545
rect 2555 2505 2595 2545
rect 2355 2205 2395 2245
rect 2955 2205 2995 2245
rect 1555 2005 1595 2045
rect 2155 2005 2195 2045
rect -45 1605 -5 1645
rect 555 1605 595 1645
rect 755 1405 795 1445
rect 1355 1405 1395 1445
rect 155 1105 195 1145
rect 1155 1105 1195 1145
rect 1755 1105 1795 1145
rect 2755 1105 2795 1145
<< metal4 >>
rect 350 2545 400 2550
rect 350 2505 355 2545
rect 395 2505 400 2545
rect 350 2500 400 2505
rect 950 2545 1000 2550
rect 950 2505 955 2545
rect 995 2505 1000 2545
rect 950 2500 1000 2505
rect 1950 2545 2000 2550
rect 1950 2505 1955 2545
rect 1995 2505 2000 2545
rect 1950 2500 2000 2505
rect 2550 2545 2600 2550
rect 2550 2505 2555 2545
rect 2595 2505 2600 2545
rect 2550 2500 2600 2505
rect 2350 2245 2400 2250
rect 2350 2205 2355 2245
rect 2395 2205 2400 2245
rect 2350 2200 2400 2205
rect 2950 2245 3000 2250
rect 2950 2205 2955 2245
rect 2995 2205 3000 2245
rect 2950 2200 3000 2205
rect 1550 2045 1600 2050
rect 1550 2005 1555 2045
rect 1595 2005 1600 2045
rect 1550 2000 1600 2005
rect 2150 2045 2200 2050
rect 2150 2005 2155 2045
rect 2195 2005 2200 2045
rect 2150 2000 2200 2005
rect -50 1645 0 1650
rect -50 1605 -45 1645
rect -5 1605 0 1645
rect -50 1600 0 1605
rect 550 1645 600 1650
rect 550 1605 555 1645
rect 595 1605 600 1645
rect 550 1600 600 1605
rect 750 1445 800 1450
rect 750 1405 755 1445
rect 795 1405 800 1445
rect 750 1400 800 1405
rect 1350 1445 1400 1450
rect 1350 1405 1355 1445
rect 1395 1405 1400 1445
rect 1350 1400 1400 1405
rect 150 1145 200 1150
rect 150 1105 155 1145
rect 195 1105 200 1145
rect 150 1100 200 1105
rect 1150 1145 1200 1150
rect 1150 1105 1155 1145
rect 1195 1105 1200 1145
rect 1150 1100 1200 1105
rect 1750 1145 1800 1150
rect 1750 1105 1755 1145
rect 1795 1105 1800 1145
rect 1750 1100 1800 1105
rect 2750 1145 2800 1150
rect 2750 1105 2755 1145
rect 2795 1105 2800 1145
rect 2750 1100 2800 1105
use inv1x  aam
timestamp 1719349823
transform 1 0 700 0 1 1050
box -100 -1150 250 2700
use inv1x  aap
timestamp 1719349823
transform 1 0 -100 0 1 1050
box -100 -1150 250 2700
use inv1x  abm
timestamp 1719349823
transform -1 0 1450 0 1 1050
box -100 -1150 250 2700
use inv1x  abp
timestamp 1719349823
transform -1 0 650 0 1 1050
box -100 -1150 250 2700
use inv1x  acm
timestamp 1719349823
transform -1 0 1050 0 1 1050
box -100 -1150 250 2700
use inv1x  acp
timestamp 1719349823
transform -1 0 250 0 1 1050
box -100 -1150 250 2700
use inv1x  adm
timestamp 1719349823
transform 1 0 1100 0 1 1050
box -100 -1150 250 2700
use inv1x  adp
timestamp 1719349823
transform 1 0 300 0 1 1050
box -100 -1150 250 2700
use inv1x  bam
timestamp 1719349823
transform 1 0 2300 0 1 1050
box -100 -1150 250 2700
use inv1x  bap
timestamp 1719349823
transform 1 0 1500 0 1 1050
box -100 -1150 250 2700
use inv1x  bbm
timestamp 1719349823
transform -1 0 3050 0 1 1050
box -100 -1150 250 2700
use inv1x  bbp
timestamp 1719349823
transform -1 0 2250 0 1 1050
box -100 -1150 250 2700
use inv1x  bcm
timestamp 1719349823
transform -1 0 2650 0 1 1050
box -100 -1150 250 2700
use inv1x  bcp
timestamp 1719349823
transform -1 0 1850 0 1 1050
box -100 -1150 250 2700
use inv1x  bdm
timestamp 1719349823
transform 1 0 2700 0 1 1050
box -100 -1150 250 2700
use inv1x  bdp
timestamp 1719349823
transform 1 0 1900 0 1 1050
box -100 -1150 250 2700
<< labels >>
rlabel metal3 -150 1600 3100 1650 0 ipa
port 1 nsew
rlabel metal3 -150 1400 3100 1450 0 ima
port 2 nsew
rlabel metal3 -150 2000 3100 2050 0 ipb
port 3 nsew
rlabel metal3 -150 2200 3100 2250 0 imb
port 4 nsew
rlabel metal3 -150 2400 3100 2650 0 op
port 5 nsew
rlabel metal3 -150 1000 3100 1250 0 om
port 6 nsew
rlabel locali -150 50 3050 100 0 bp
port 7 nsew
rlabel locali -150 950 3100 1000 0 bn
port 8 nsew
rlabel metal3 -150 2700 3100 2750 0 vss
port 10 nsew
rlabel locali -200 -100 3150 -50 0 vsub
port 11 nsew
rlabel locali -100 950 -50 1000 0 bn
<< end >>
