magic
tech sky130A
timestamp 1725883591
<< dnwell >>
rect 1595 895 2955 2955
<< nwell >>
rect 1550 2850 3000 3750
rect 1550 1000 1700 2850
rect 2850 1000 3000 2850
rect 1550 100 3000 1000
<< pwell >>
rect 1850 2800 2700 2850
rect 1750 2750 2800 2800
rect 1750 1100 1800 2750
rect 1850 2000 2700 2750
rect 1850 1850 2050 2000
rect 2100 1850 2450 2000
rect 2500 1850 2700 2000
rect 1850 1100 2700 1850
rect 2750 1100 2800 2750
rect 1750 1050 2800 1100
rect 1850 1000 2700 1050
<< pmoslvt >>
rect 1900 3100 1950 3600
rect 2000 3100 2050 3600
rect 2100 3100 2150 3600
rect 2200 3100 2250 3600
rect 2300 3100 2350 3600
rect 2400 3100 2450 3600
rect 2500 3100 2550 3600
rect 2600 3100 2650 3600
rect 1900 250 1950 750
rect 2000 250 2050 750
rect 2100 250 2150 750
rect 2200 250 2250 750
rect 2300 250 2350 750
rect 2400 250 2450 750
rect 2500 250 2550 750
rect 2600 250 2650 750
<< nmoslvt >>
rect 1900 2000 1950 2700
rect 2000 2000 2050 2700
rect 2100 2000 2150 2700
rect 2200 2000 2250 2700
rect 2300 2000 2350 2700
rect 2400 2000 2450 2700
rect 2500 2000 2550 2700
rect 2600 2000 2650 2700
rect 1900 1150 1950 1850
rect 2000 1150 2050 1850
rect 2100 1150 2150 1850
rect 2200 1150 2250 1850
rect 2300 1150 2350 1850
rect 2400 1150 2450 1850
rect 2500 1150 2550 1850
rect 2600 1150 2650 1850
<< ndiff >>
rect 1850 2685 1900 2700
rect 1850 2665 1865 2685
rect 1885 2665 1900 2685
rect 1850 2635 1900 2665
rect 1850 2615 1865 2635
rect 1885 2615 1900 2635
rect 1850 2585 1900 2615
rect 1850 2565 1865 2585
rect 1885 2565 1900 2585
rect 1850 2535 1900 2565
rect 1850 2515 1865 2535
rect 1885 2515 1900 2535
rect 1850 2485 1900 2515
rect 1850 2465 1865 2485
rect 1885 2465 1900 2485
rect 1850 2435 1900 2465
rect 1850 2415 1865 2435
rect 1885 2415 1900 2435
rect 1850 2385 1900 2415
rect 1850 2365 1865 2385
rect 1885 2365 1900 2385
rect 1850 2335 1900 2365
rect 1850 2315 1865 2335
rect 1885 2315 1900 2335
rect 1850 2285 1900 2315
rect 1850 2265 1865 2285
rect 1885 2265 1900 2285
rect 1850 2235 1900 2265
rect 1850 2215 1865 2235
rect 1885 2215 1900 2235
rect 1850 2185 1900 2215
rect 1850 2165 1865 2185
rect 1885 2165 1900 2185
rect 1850 2135 1900 2165
rect 1850 2115 1865 2135
rect 1885 2115 1900 2135
rect 1850 2085 1900 2115
rect 1850 2065 1865 2085
rect 1885 2065 1900 2085
rect 1850 2035 1900 2065
rect 1850 2015 1865 2035
rect 1885 2015 1900 2035
rect 1850 2000 1900 2015
rect 1950 2000 2000 2700
rect 2050 2685 2100 2700
rect 2050 2665 2065 2685
rect 2085 2665 2100 2685
rect 2050 2635 2100 2665
rect 2050 2615 2065 2635
rect 2085 2615 2100 2635
rect 2050 2585 2100 2615
rect 2050 2565 2065 2585
rect 2085 2565 2100 2585
rect 2050 2535 2100 2565
rect 2050 2515 2065 2535
rect 2085 2515 2100 2535
rect 2050 2485 2100 2515
rect 2050 2465 2065 2485
rect 2085 2465 2100 2485
rect 2050 2435 2100 2465
rect 2050 2415 2065 2435
rect 2085 2415 2100 2435
rect 2050 2385 2100 2415
rect 2050 2365 2065 2385
rect 2085 2365 2100 2385
rect 2050 2335 2100 2365
rect 2050 2315 2065 2335
rect 2085 2315 2100 2335
rect 2050 2285 2100 2315
rect 2050 2265 2065 2285
rect 2085 2265 2100 2285
rect 2050 2235 2100 2265
rect 2050 2215 2065 2235
rect 2085 2215 2100 2235
rect 2050 2185 2100 2215
rect 2050 2165 2065 2185
rect 2085 2165 2100 2185
rect 2050 2135 2100 2165
rect 2050 2115 2065 2135
rect 2085 2115 2100 2135
rect 2050 2085 2100 2115
rect 2050 2065 2065 2085
rect 2085 2065 2100 2085
rect 2050 2035 2100 2065
rect 2050 2015 2065 2035
rect 2085 2015 2100 2035
rect 2050 2000 2100 2015
rect 2150 2000 2200 2700
rect 2250 2685 2300 2700
rect 2250 2665 2265 2685
rect 2285 2665 2300 2685
rect 2250 2635 2300 2665
rect 2250 2615 2265 2635
rect 2285 2615 2300 2635
rect 2250 2585 2300 2615
rect 2250 2565 2265 2585
rect 2285 2565 2300 2585
rect 2250 2535 2300 2565
rect 2250 2515 2265 2535
rect 2285 2515 2300 2535
rect 2250 2485 2300 2515
rect 2250 2465 2265 2485
rect 2285 2465 2300 2485
rect 2250 2435 2300 2465
rect 2250 2415 2265 2435
rect 2285 2415 2300 2435
rect 2250 2385 2300 2415
rect 2250 2365 2265 2385
rect 2285 2365 2300 2385
rect 2250 2335 2300 2365
rect 2250 2315 2265 2335
rect 2285 2315 2300 2335
rect 2250 2285 2300 2315
rect 2250 2265 2265 2285
rect 2285 2265 2300 2285
rect 2250 2235 2300 2265
rect 2250 2215 2265 2235
rect 2285 2215 2300 2235
rect 2250 2185 2300 2215
rect 2250 2165 2265 2185
rect 2285 2165 2300 2185
rect 2250 2135 2300 2165
rect 2250 2115 2265 2135
rect 2285 2115 2300 2135
rect 2250 2085 2300 2115
rect 2250 2065 2265 2085
rect 2285 2065 2300 2085
rect 2250 2035 2300 2065
rect 2250 2015 2265 2035
rect 2285 2015 2300 2035
rect 2250 2000 2300 2015
rect 2350 2000 2400 2700
rect 2450 2685 2500 2700
rect 2450 2665 2465 2685
rect 2485 2665 2500 2685
rect 2450 2635 2500 2665
rect 2450 2615 2465 2635
rect 2485 2615 2500 2635
rect 2450 2585 2500 2615
rect 2450 2565 2465 2585
rect 2485 2565 2500 2585
rect 2450 2535 2500 2565
rect 2450 2515 2465 2535
rect 2485 2515 2500 2535
rect 2450 2485 2500 2515
rect 2450 2465 2465 2485
rect 2485 2465 2500 2485
rect 2450 2435 2500 2465
rect 2450 2415 2465 2435
rect 2485 2415 2500 2435
rect 2450 2385 2500 2415
rect 2450 2365 2465 2385
rect 2485 2365 2500 2385
rect 2450 2335 2500 2365
rect 2450 2315 2465 2335
rect 2485 2315 2500 2335
rect 2450 2285 2500 2315
rect 2450 2265 2465 2285
rect 2485 2265 2500 2285
rect 2450 2235 2500 2265
rect 2450 2215 2465 2235
rect 2485 2215 2500 2235
rect 2450 2185 2500 2215
rect 2450 2165 2465 2185
rect 2485 2165 2500 2185
rect 2450 2135 2500 2165
rect 2450 2115 2465 2135
rect 2485 2115 2500 2135
rect 2450 2085 2500 2115
rect 2450 2065 2465 2085
rect 2485 2065 2500 2085
rect 2450 2035 2500 2065
rect 2450 2015 2465 2035
rect 2485 2015 2500 2035
rect 2450 2000 2500 2015
rect 2550 2000 2600 2700
rect 2650 2685 2700 2700
rect 2650 2665 2665 2685
rect 2685 2665 2700 2685
rect 2650 2635 2700 2665
rect 2650 2615 2665 2635
rect 2685 2615 2700 2635
rect 2650 2585 2700 2615
rect 2650 2565 2665 2585
rect 2685 2565 2700 2585
rect 2650 2535 2700 2565
rect 2650 2515 2665 2535
rect 2685 2515 2700 2535
rect 2650 2485 2700 2515
rect 2650 2465 2665 2485
rect 2685 2465 2700 2485
rect 2650 2435 2700 2465
rect 2650 2415 2665 2435
rect 2685 2415 2700 2435
rect 2650 2385 2700 2415
rect 2650 2365 2665 2385
rect 2685 2365 2700 2385
rect 2650 2335 2700 2365
rect 2650 2315 2665 2335
rect 2685 2315 2700 2335
rect 2650 2285 2700 2315
rect 2650 2265 2665 2285
rect 2685 2265 2700 2285
rect 2650 2235 2700 2265
rect 2650 2215 2665 2235
rect 2685 2215 2700 2235
rect 2650 2185 2700 2215
rect 2650 2165 2665 2185
rect 2685 2165 2700 2185
rect 2650 2135 2700 2165
rect 2650 2115 2665 2135
rect 2685 2115 2700 2135
rect 2650 2085 2700 2115
rect 2650 2065 2665 2085
rect 2685 2065 2700 2085
rect 2650 2035 2700 2065
rect 2650 2015 2665 2035
rect 2685 2015 2700 2035
rect 2650 2000 2700 2015
rect 1850 1835 1900 1850
rect 1850 1815 1865 1835
rect 1885 1815 1900 1835
rect 1850 1785 1900 1815
rect 1850 1765 1865 1785
rect 1885 1765 1900 1785
rect 1850 1735 1900 1765
rect 1850 1715 1865 1735
rect 1885 1715 1900 1735
rect 1850 1685 1900 1715
rect 1850 1665 1865 1685
rect 1885 1665 1900 1685
rect 1850 1635 1900 1665
rect 1850 1615 1865 1635
rect 1885 1615 1900 1635
rect 1850 1585 1900 1615
rect 1850 1565 1865 1585
rect 1885 1565 1900 1585
rect 1850 1535 1900 1565
rect 1850 1515 1865 1535
rect 1885 1515 1900 1535
rect 1850 1485 1900 1515
rect 1850 1465 1865 1485
rect 1885 1465 1900 1485
rect 1850 1435 1900 1465
rect 1850 1415 1865 1435
rect 1885 1415 1900 1435
rect 1850 1385 1900 1415
rect 1850 1365 1865 1385
rect 1885 1365 1900 1385
rect 1850 1335 1900 1365
rect 1850 1315 1865 1335
rect 1885 1315 1900 1335
rect 1850 1285 1900 1315
rect 1850 1265 1865 1285
rect 1885 1265 1900 1285
rect 1850 1235 1900 1265
rect 1850 1215 1865 1235
rect 1885 1215 1900 1235
rect 1850 1185 1900 1215
rect 1850 1165 1865 1185
rect 1885 1165 1900 1185
rect 1850 1150 1900 1165
rect 1950 1150 2000 1850
rect 2050 1835 2100 1850
rect 2050 1815 2065 1835
rect 2085 1815 2100 1835
rect 2050 1785 2100 1815
rect 2050 1765 2065 1785
rect 2085 1765 2100 1785
rect 2050 1735 2100 1765
rect 2050 1715 2065 1735
rect 2085 1715 2100 1735
rect 2050 1685 2100 1715
rect 2050 1665 2065 1685
rect 2085 1665 2100 1685
rect 2050 1635 2100 1665
rect 2050 1615 2065 1635
rect 2085 1615 2100 1635
rect 2050 1585 2100 1615
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1150 2100 1165
rect 2150 1150 2200 1850
rect 2250 1835 2300 1850
rect 2250 1815 2265 1835
rect 2285 1815 2300 1835
rect 2250 1785 2300 1815
rect 2250 1765 2265 1785
rect 2285 1765 2300 1785
rect 2250 1735 2300 1765
rect 2250 1715 2265 1735
rect 2285 1715 2300 1735
rect 2250 1685 2300 1715
rect 2250 1665 2265 1685
rect 2285 1665 2300 1685
rect 2250 1635 2300 1665
rect 2250 1615 2265 1635
rect 2285 1615 2300 1635
rect 2250 1585 2300 1615
rect 2250 1565 2265 1585
rect 2285 1565 2300 1585
rect 2250 1535 2300 1565
rect 2250 1515 2265 1535
rect 2285 1515 2300 1535
rect 2250 1485 2300 1515
rect 2250 1465 2265 1485
rect 2285 1465 2300 1485
rect 2250 1435 2300 1465
rect 2250 1415 2265 1435
rect 2285 1415 2300 1435
rect 2250 1385 2300 1415
rect 2250 1365 2265 1385
rect 2285 1365 2300 1385
rect 2250 1335 2300 1365
rect 2250 1315 2265 1335
rect 2285 1315 2300 1335
rect 2250 1285 2300 1315
rect 2250 1265 2265 1285
rect 2285 1265 2300 1285
rect 2250 1235 2300 1265
rect 2250 1215 2265 1235
rect 2285 1215 2300 1235
rect 2250 1185 2300 1215
rect 2250 1165 2265 1185
rect 2285 1165 2300 1185
rect 2250 1150 2300 1165
rect 2350 1150 2400 1850
rect 2450 1835 2500 1850
rect 2450 1815 2465 1835
rect 2485 1815 2500 1835
rect 2450 1785 2500 1815
rect 2450 1765 2465 1785
rect 2485 1765 2500 1785
rect 2450 1735 2500 1765
rect 2450 1715 2465 1735
rect 2485 1715 2500 1735
rect 2450 1685 2500 1715
rect 2450 1665 2465 1685
rect 2485 1665 2500 1685
rect 2450 1635 2500 1665
rect 2450 1615 2465 1635
rect 2485 1615 2500 1635
rect 2450 1585 2500 1615
rect 2450 1565 2465 1585
rect 2485 1565 2500 1585
rect 2450 1535 2500 1565
rect 2450 1515 2465 1535
rect 2485 1515 2500 1535
rect 2450 1485 2500 1515
rect 2450 1465 2465 1485
rect 2485 1465 2500 1485
rect 2450 1435 2500 1465
rect 2450 1415 2465 1435
rect 2485 1415 2500 1435
rect 2450 1385 2500 1415
rect 2450 1365 2465 1385
rect 2485 1365 2500 1385
rect 2450 1335 2500 1365
rect 2450 1315 2465 1335
rect 2485 1315 2500 1335
rect 2450 1285 2500 1315
rect 2450 1265 2465 1285
rect 2485 1265 2500 1285
rect 2450 1235 2500 1265
rect 2450 1215 2465 1235
rect 2485 1215 2500 1235
rect 2450 1185 2500 1215
rect 2450 1165 2465 1185
rect 2485 1165 2500 1185
rect 2450 1150 2500 1165
rect 2550 1150 2600 1850
rect 2650 1835 2700 1850
rect 2650 1815 2665 1835
rect 2685 1815 2700 1835
rect 2650 1785 2700 1815
rect 2650 1765 2665 1785
rect 2685 1765 2700 1785
rect 2650 1735 2700 1765
rect 2650 1715 2665 1735
rect 2685 1715 2700 1735
rect 2650 1685 2700 1715
rect 2650 1665 2665 1685
rect 2685 1665 2700 1685
rect 2650 1635 2700 1665
rect 2650 1615 2665 1635
rect 2685 1615 2700 1635
rect 2650 1585 2700 1615
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1150 2700 1165
<< pdiff >>
rect 1850 3585 1900 3600
rect 1850 3565 1865 3585
rect 1885 3565 1900 3585
rect 1850 3535 1900 3565
rect 1850 3515 1865 3535
rect 1885 3515 1900 3535
rect 1850 3485 1900 3515
rect 1850 3465 1865 3485
rect 1885 3465 1900 3485
rect 1850 3435 1900 3465
rect 1850 3415 1865 3435
rect 1885 3415 1900 3435
rect 1850 3385 1900 3415
rect 1850 3365 1865 3385
rect 1885 3365 1900 3385
rect 1850 3335 1900 3365
rect 1850 3315 1865 3335
rect 1885 3315 1900 3335
rect 1850 3285 1900 3315
rect 1850 3265 1865 3285
rect 1885 3265 1900 3285
rect 1850 3235 1900 3265
rect 1850 3215 1865 3235
rect 1885 3215 1900 3235
rect 1850 3185 1900 3215
rect 1850 3165 1865 3185
rect 1885 3165 1900 3185
rect 1850 3135 1900 3165
rect 1850 3115 1865 3135
rect 1885 3115 1900 3135
rect 1850 3100 1900 3115
rect 1950 3585 2000 3600
rect 1950 3565 1965 3585
rect 1985 3565 2000 3585
rect 1950 3535 2000 3565
rect 1950 3515 1965 3535
rect 1985 3515 2000 3535
rect 1950 3485 2000 3515
rect 1950 3465 1965 3485
rect 1985 3465 2000 3485
rect 1950 3435 2000 3465
rect 1950 3415 1965 3435
rect 1985 3415 2000 3435
rect 1950 3385 2000 3415
rect 1950 3365 1965 3385
rect 1985 3365 2000 3385
rect 1950 3335 2000 3365
rect 1950 3315 1965 3335
rect 1985 3315 2000 3335
rect 1950 3285 2000 3315
rect 1950 3265 1965 3285
rect 1985 3265 2000 3285
rect 1950 3235 2000 3265
rect 1950 3215 1965 3235
rect 1985 3215 2000 3235
rect 1950 3185 2000 3215
rect 1950 3165 1965 3185
rect 1985 3165 2000 3185
rect 1950 3135 2000 3165
rect 1950 3115 1965 3135
rect 1985 3115 2000 3135
rect 1950 3100 2000 3115
rect 2050 3585 2100 3600
rect 2050 3565 2065 3585
rect 2085 3565 2100 3585
rect 2050 3535 2100 3565
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3285 2100 3315
rect 2050 3265 2065 3285
rect 2085 3265 2100 3285
rect 2050 3235 2100 3265
rect 2050 3215 2065 3235
rect 2085 3215 2100 3235
rect 2050 3185 2100 3215
rect 2050 3165 2065 3185
rect 2085 3165 2100 3185
rect 2050 3135 2100 3165
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3100 2100 3115
rect 2150 3585 2200 3600
rect 2150 3565 2165 3585
rect 2185 3565 2200 3585
rect 2150 3535 2200 3565
rect 2150 3515 2165 3535
rect 2185 3515 2200 3535
rect 2150 3485 2200 3515
rect 2150 3465 2165 3485
rect 2185 3465 2200 3485
rect 2150 3435 2200 3465
rect 2150 3415 2165 3435
rect 2185 3415 2200 3435
rect 2150 3385 2200 3415
rect 2150 3365 2165 3385
rect 2185 3365 2200 3385
rect 2150 3335 2200 3365
rect 2150 3315 2165 3335
rect 2185 3315 2200 3335
rect 2150 3285 2200 3315
rect 2150 3265 2165 3285
rect 2185 3265 2200 3285
rect 2150 3235 2200 3265
rect 2150 3215 2165 3235
rect 2185 3215 2200 3235
rect 2150 3185 2200 3215
rect 2150 3165 2165 3185
rect 2185 3165 2200 3185
rect 2150 3135 2200 3165
rect 2150 3115 2165 3135
rect 2185 3115 2200 3135
rect 2150 3100 2200 3115
rect 2250 3585 2300 3600
rect 2250 3565 2265 3585
rect 2285 3565 2300 3585
rect 2250 3535 2300 3565
rect 2250 3515 2265 3535
rect 2285 3515 2300 3535
rect 2250 3485 2300 3515
rect 2250 3465 2265 3485
rect 2285 3465 2300 3485
rect 2250 3435 2300 3465
rect 2250 3415 2265 3435
rect 2285 3415 2300 3435
rect 2250 3385 2300 3415
rect 2250 3365 2265 3385
rect 2285 3365 2300 3385
rect 2250 3335 2300 3365
rect 2250 3315 2265 3335
rect 2285 3315 2300 3335
rect 2250 3285 2300 3315
rect 2250 3265 2265 3285
rect 2285 3265 2300 3285
rect 2250 3235 2300 3265
rect 2250 3215 2265 3235
rect 2285 3215 2300 3235
rect 2250 3185 2300 3215
rect 2250 3165 2265 3185
rect 2285 3165 2300 3185
rect 2250 3135 2300 3165
rect 2250 3115 2265 3135
rect 2285 3115 2300 3135
rect 2250 3100 2300 3115
rect 2350 3585 2400 3600
rect 2350 3565 2365 3585
rect 2385 3565 2400 3585
rect 2350 3535 2400 3565
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3285 2400 3315
rect 2350 3265 2365 3285
rect 2385 3265 2400 3285
rect 2350 3235 2400 3265
rect 2350 3215 2365 3235
rect 2385 3215 2400 3235
rect 2350 3185 2400 3215
rect 2350 3165 2365 3185
rect 2385 3165 2400 3185
rect 2350 3135 2400 3165
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3100 2400 3115
rect 2450 3585 2500 3600
rect 2450 3565 2465 3585
rect 2485 3565 2500 3585
rect 2450 3535 2500 3565
rect 2450 3515 2465 3535
rect 2485 3515 2500 3535
rect 2450 3485 2500 3515
rect 2450 3465 2465 3485
rect 2485 3465 2500 3485
rect 2450 3435 2500 3465
rect 2450 3415 2465 3435
rect 2485 3415 2500 3435
rect 2450 3385 2500 3415
rect 2450 3365 2465 3385
rect 2485 3365 2500 3385
rect 2450 3335 2500 3365
rect 2450 3315 2465 3335
rect 2485 3315 2500 3335
rect 2450 3285 2500 3315
rect 2450 3265 2465 3285
rect 2485 3265 2500 3285
rect 2450 3235 2500 3265
rect 2450 3215 2465 3235
rect 2485 3215 2500 3235
rect 2450 3185 2500 3215
rect 2450 3165 2465 3185
rect 2485 3165 2500 3185
rect 2450 3135 2500 3165
rect 2450 3115 2465 3135
rect 2485 3115 2500 3135
rect 2450 3100 2500 3115
rect 2550 3585 2600 3600
rect 2550 3565 2565 3585
rect 2585 3565 2600 3585
rect 2550 3535 2600 3565
rect 2550 3515 2565 3535
rect 2585 3515 2600 3535
rect 2550 3485 2600 3515
rect 2550 3465 2565 3485
rect 2585 3465 2600 3485
rect 2550 3435 2600 3465
rect 2550 3415 2565 3435
rect 2585 3415 2600 3435
rect 2550 3385 2600 3415
rect 2550 3365 2565 3385
rect 2585 3365 2600 3385
rect 2550 3335 2600 3365
rect 2550 3315 2565 3335
rect 2585 3315 2600 3335
rect 2550 3285 2600 3315
rect 2550 3265 2565 3285
rect 2585 3265 2600 3285
rect 2550 3235 2600 3265
rect 2550 3215 2565 3235
rect 2585 3215 2600 3235
rect 2550 3185 2600 3215
rect 2550 3165 2565 3185
rect 2585 3165 2600 3185
rect 2550 3135 2600 3165
rect 2550 3115 2565 3135
rect 2585 3115 2600 3135
rect 2550 3100 2600 3115
rect 2650 3585 2700 3600
rect 2650 3565 2665 3585
rect 2685 3565 2700 3585
rect 2650 3535 2700 3565
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3285 2700 3315
rect 2650 3265 2665 3285
rect 2685 3265 2700 3285
rect 2650 3235 2700 3265
rect 2650 3215 2665 3235
rect 2685 3215 2700 3235
rect 2650 3185 2700 3215
rect 2650 3165 2665 3185
rect 2685 3165 2700 3185
rect 2650 3135 2700 3165
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3100 2700 3115
rect 1850 735 1900 750
rect 1850 715 1865 735
rect 1885 715 1900 735
rect 1850 685 1900 715
rect 1850 665 1865 685
rect 1885 665 1900 685
rect 1850 635 1900 665
rect 1850 615 1865 635
rect 1885 615 1900 635
rect 1850 585 1900 615
rect 1850 565 1865 585
rect 1885 565 1900 585
rect 1850 535 1900 565
rect 1850 515 1865 535
rect 1885 515 1900 535
rect 1850 485 1900 515
rect 1850 465 1865 485
rect 1885 465 1900 485
rect 1850 435 1900 465
rect 1850 415 1865 435
rect 1885 415 1900 435
rect 1850 385 1900 415
rect 1850 365 1865 385
rect 1885 365 1900 385
rect 1850 335 1900 365
rect 1850 315 1865 335
rect 1885 315 1900 335
rect 1850 285 1900 315
rect 1850 265 1865 285
rect 1885 265 1900 285
rect 1850 250 1900 265
rect 1950 735 2000 750
rect 1950 715 1965 735
rect 1985 715 2000 735
rect 1950 685 2000 715
rect 1950 665 1965 685
rect 1985 665 2000 685
rect 1950 635 2000 665
rect 1950 615 1965 635
rect 1985 615 2000 635
rect 1950 585 2000 615
rect 1950 565 1965 585
rect 1985 565 2000 585
rect 1950 535 2000 565
rect 1950 515 1965 535
rect 1985 515 2000 535
rect 1950 485 2000 515
rect 1950 465 1965 485
rect 1985 465 2000 485
rect 1950 435 2000 465
rect 1950 415 1965 435
rect 1985 415 2000 435
rect 1950 385 2000 415
rect 1950 365 1965 385
rect 1985 365 2000 385
rect 1950 335 2000 365
rect 1950 315 1965 335
rect 1985 315 2000 335
rect 1950 285 2000 315
rect 1950 265 1965 285
rect 1985 265 2000 285
rect 1950 250 2000 265
rect 2050 735 2100 750
rect 2050 715 2065 735
rect 2085 715 2100 735
rect 2050 685 2100 715
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 2050 635 2100 665
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 250 2100 265
rect 2150 735 2200 750
rect 2150 715 2165 735
rect 2185 715 2200 735
rect 2150 685 2200 715
rect 2150 665 2165 685
rect 2185 665 2200 685
rect 2150 635 2200 665
rect 2150 615 2165 635
rect 2185 615 2200 635
rect 2150 585 2200 615
rect 2150 565 2165 585
rect 2185 565 2200 585
rect 2150 535 2200 565
rect 2150 515 2165 535
rect 2185 515 2200 535
rect 2150 485 2200 515
rect 2150 465 2165 485
rect 2185 465 2200 485
rect 2150 435 2200 465
rect 2150 415 2165 435
rect 2185 415 2200 435
rect 2150 385 2200 415
rect 2150 365 2165 385
rect 2185 365 2200 385
rect 2150 335 2200 365
rect 2150 315 2165 335
rect 2185 315 2200 335
rect 2150 285 2200 315
rect 2150 265 2165 285
rect 2185 265 2200 285
rect 2150 250 2200 265
rect 2250 735 2300 750
rect 2250 715 2265 735
rect 2285 715 2300 735
rect 2250 685 2300 715
rect 2250 665 2265 685
rect 2285 665 2300 685
rect 2250 635 2300 665
rect 2250 615 2265 635
rect 2285 615 2300 635
rect 2250 585 2300 615
rect 2250 565 2265 585
rect 2285 565 2300 585
rect 2250 535 2300 565
rect 2250 515 2265 535
rect 2285 515 2300 535
rect 2250 485 2300 515
rect 2250 465 2265 485
rect 2285 465 2300 485
rect 2250 435 2300 465
rect 2250 415 2265 435
rect 2285 415 2300 435
rect 2250 385 2300 415
rect 2250 365 2265 385
rect 2285 365 2300 385
rect 2250 335 2300 365
rect 2250 315 2265 335
rect 2285 315 2300 335
rect 2250 285 2300 315
rect 2250 265 2265 285
rect 2285 265 2300 285
rect 2250 250 2300 265
rect 2350 735 2400 750
rect 2350 715 2365 735
rect 2385 715 2400 735
rect 2350 685 2400 715
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 250 2400 265
rect 2450 735 2500 750
rect 2450 715 2465 735
rect 2485 715 2500 735
rect 2450 685 2500 715
rect 2450 665 2465 685
rect 2485 665 2500 685
rect 2450 635 2500 665
rect 2450 615 2465 635
rect 2485 615 2500 635
rect 2450 585 2500 615
rect 2450 565 2465 585
rect 2485 565 2500 585
rect 2450 535 2500 565
rect 2450 515 2465 535
rect 2485 515 2500 535
rect 2450 485 2500 515
rect 2450 465 2465 485
rect 2485 465 2500 485
rect 2450 435 2500 465
rect 2450 415 2465 435
rect 2485 415 2500 435
rect 2450 385 2500 415
rect 2450 365 2465 385
rect 2485 365 2500 385
rect 2450 335 2500 365
rect 2450 315 2465 335
rect 2485 315 2500 335
rect 2450 285 2500 315
rect 2450 265 2465 285
rect 2485 265 2500 285
rect 2450 250 2500 265
rect 2550 735 2600 750
rect 2550 715 2565 735
rect 2585 715 2600 735
rect 2550 685 2600 715
rect 2550 665 2565 685
rect 2585 665 2600 685
rect 2550 635 2600 665
rect 2550 615 2565 635
rect 2585 615 2600 635
rect 2550 585 2600 615
rect 2550 565 2565 585
rect 2585 565 2600 585
rect 2550 535 2600 565
rect 2550 515 2565 535
rect 2585 515 2600 535
rect 2550 485 2600 515
rect 2550 465 2565 485
rect 2585 465 2600 485
rect 2550 435 2600 465
rect 2550 415 2565 435
rect 2585 415 2600 435
rect 2550 385 2600 415
rect 2550 365 2565 385
rect 2585 365 2600 385
rect 2550 335 2600 365
rect 2550 315 2565 335
rect 2585 315 2600 335
rect 2550 285 2600 315
rect 2550 265 2565 285
rect 2585 265 2600 285
rect 2550 250 2600 265
rect 2650 735 2700 750
rect 2650 715 2665 735
rect 2685 715 2700 735
rect 2650 685 2700 715
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 635 2700 665
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 250 2700 265
<< ndiffc >>
rect 1865 2665 1885 2685
rect 1865 2615 1885 2635
rect 1865 2565 1885 2585
rect 1865 2515 1885 2535
rect 1865 2465 1885 2485
rect 1865 2415 1885 2435
rect 1865 2365 1885 2385
rect 1865 2315 1885 2335
rect 1865 2265 1885 2285
rect 1865 2215 1885 2235
rect 1865 2165 1885 2185
rect 1865 2115 1885 2135
rect 1865 2065 1885 2085
rect 1865 2015 1885 2035
rect 2065 2665 2085 2685
rect 2065 2615 2085 2635
rect 2065 2565 2085 2585
rect 2065 2515 2085 2535
rect 2065 2465 2085 2485
rect 2065 2415 2085 2435
rect 2065 2365 2085 2385
rect 2065 2315 2085 2335
rect 2065 2265 2085 2285
rect 2065 2215 2085 2235
rect 2065 2165 2085 2185
rect 2065 2115 2085 2135
rect 2065 2065 2085 2085
rect 2065 2015 2085 2035
rect 2265 2665 2285 2685
rect 2265 2615 2285 2635
rect 2265 2565 2285 2585
rect 2265 2515 2285 2535
rect 2265 2465 2285 2485
rect 2265 2415 2285 2435
rect 2265 2365 2285 2385
rect 2265 2315 2285 2335
rect 2265 2265 2285 2285
rect 2265 2215 2285 2235
rect 2265 2165 2285 2185
rect 2265 2115 2285 2135
rect 2265 2065 2285 2085
rect 2265 2015 2285 2035
rect 2465 2665 2485 2685
rect 2465 2615 2485 2635
rect 2465 2565 2485 2585
rect 2465 2515 2485 2535
rect 2465 2465 2485 2485
rect 2465 2415 2485 2435
rect 2465 2365 2485 2385
rect 2465 2315 2485 2335
rect 2465 2265 2485 2285
rect 2465 2215 2485 2235
rect 2465 2165 2485 2185
rect 2465 2115 2485 2135
rect 2465 2065 2485 2085
rect 2465 2015 2485 2035
rect 2665 2665 2685 2685
rect 2665 2615 2685 2635
rect 2665 2565 2685 2585
rect 2665 2515 2685 2535
rect 2665 2465 2685 2485
rect 2665 2415 2685 2435
rect 2665 2365 2685 2385
rect 2665 2315 2685 2335
rect 2665 2265 2685 2285
rect 2665 2215 2685 2235
rect 2665 2165 2685 2185
rect 2665 2115 2685 2135
rect 2665 2065 2685 2085
rect 2665 2015 2685 2035
rect 1865 1815 1885 1835
rect 1865 1765 1885 1785
rect 1865 1715 1885 1735
rect 1865 1665 1885 1685
rect 1865 1615 1885 1635
rect 1865 1565 1885 1585
rect 1865 1515 1885 1535
rect 1865 1465 1885 1485
rect 1865 1415 1885 1435
rect 1865 1365 1885 1385
rect 1865 1315 1885 1335
rect 1865 1265 1885 1285
rect 1865 1215 1885 1235
rect 1865 1165 1885 1185
rect 2065 1815 2085 1835
rect 2065 1765 2085 1785
rect 2065 1715 2085 1735
rect 2065 1665 2085 1685
rect 2065 1615 2085 1635
rect 2065 1565 2085 1585
rect 2065 1515 2085 1535
rect 2065 1465 2085 1485
rect 2065 1415 2085 1435
rect 2065 1365 2085 1385
rect 2065 1315 2085 1335
rect 2065 1265 2085 1285
rect 2065 1215 2085 1235
rect 2065 1165 2085 1185
rect 2265 1815 2285 1835
rect 2265 1765 2285 1785
rect 2265 1715 2285 1735
rect 2265 1665 2285 1685
rect 2265 1615 2285 1635
rect 2265 1565 2285 1585
rect 2265 1515 2285 1535
rect 2265 1465 2285 1485
rect 2265 1415 2285 1435
rect 2265 1365 2285 1385
rect 2265 1315 2285 1335
rect 2265 1265 2285 1285
rect 2265 1215 2285 1235
rect 2265 1165 2285 1185
rect 2465 1815 2485 1835
rect 2465 1765 2485 1785
rect 2465 1715 2485 1735
rect 2465 1665 2485 1685
rect 2465 1615 2485 1635
rect 2465 1565 2485 1585
rect 2465 1515 2485 1535
rect 2465 1465 2485 1485
rect 2465 1415 2485 1435
rect 2465 1365 2485 1385
rect 2465 1315 2485 1335
rect 2465 1265 2485 1285
rect 2465 1215 2485 1235
rect 2465 1165 2485 1185
rect 2665 1815 2685 1835
rect 2665 1765 2685 1785
rect 2665 1715 2685 1735
rect 2665 1665 2685 1685
rect 2665 1615 2685 1635
rect 2665 1565 2685 1585
rect 2665 1515 2685 1535
rect 2665 1465 2685 1485
rect 2665 1415 2685 1435
rect 2665 1365 2685 1385
rect 2665 1315 2685 1335
rect 2665 1265 2685 1285
rect 2665 1215 2685 1235
rect 2665 1165 2685 1185
<< pdiffc >>
rect 1865 3565 1885 3585
rect 1865 3515 1885 3535
rect 1865 3465 1885 3485
rect 1865 3415 1885 3435
rect 1865 3365 1885 3385
rect 1865 3315 1885 3335
rect 1865 3265 1885 3285
rect 1865 3215 1885 3235
rect 1865 3165 1885 3185
rect 1865 3115 1885 3135
rect 1965 3565 1985 3585
rect 1965 3515 1985 3535
rect 1965 3465 1985 3485
rect 1965 3415 1985 3435
rect 1965 3365 1985 3385
rect 1965 3315 1985 3335
rect 1965 3265 1985 3285
rect 1965 3215 1985 3235
rect 1965 3165 1985 3185
rect 1965 3115 1985 3135
rect 2065 3565 2085 3585
rect 2065 3515 2085 3535
rect 2065 3465 2085 3485
rect 2065 3415 2085 3435
rect 2065 3365 2085 3385
rect 2065 3315 2085 3335
rect 2065 3265 2085 3285
rect 2065 3215 2085 3235
rect 2065 3165 2085 3185
rect 2065 3115 2085 3135
rect 2165 3565 2185 3585
rect 2165 3515 2185 3535
rect 2165 3465 2185 3485
rect 2165 3415 2185 3435
rect 2165 3365 2185 3385
rect 2165 3315 2185 3335
rect 2165 3265 2185 3285
rect 2165 3215 2185 3235
rect 2165 3165 2185 3185
rect 2165 3115 2185 3135
rect 2265 3565 2285 3585
rect 2265 3515 2285 3535
rect 2265 3465 2285 3485
rect 2265 3415 2285 3435
rect 2265 3365 2285 3385
rect 2265 3315 2285 3335
rect 2265 3265 2285 3285
rect 2265 3215 2285 3235
rect 2265 3165 2285 3185
rect 2265 3115 2285 3135
rect 2365 3565 2385 3585
rect 2365 3515 2385 3535
rect 2365 3465 2385 3485
rect 2365 3415 2385 3435
rect 2365 3365 2385 3385
rect 2365 3315 2385 3335
rect 2365 3265 2385 3285
rect 2365 3215 2385 3235
rect 2365 3165 2385 3185
rect 2365 3115 2385 3135
rect 2465 3565 2485 3585
rect 2465 3515 2485 3535
rect 2465 3465 2485 3485
rect 2465 3415 2485 3435
rect 2465 3365 2485 3385
rect 2465 3315 2485 3335
rect 2465 3265 2485 3285
rect 2465 3215 2485 3235
rect 2465 3165 2485 3185
rect 2465 3115 2485 3135
rect 2565 3565 2585 3585
rect 2565 3515 2585 3535
rect 2565 3465 2585 3485
rect 2565 3415 2585 3435
rect 2565 3365 2585 3385
rect 2565 3315 2585 3335
rect 2565 3265 2585 3285
rect 2565 3215 2585 3235
rect 2565 3165 2585 3185
rect 2565 3115 2585 3135
rect 2665 3565 2685 3585
rect 2665 3515 2685 3535
rect 2665 3465 2685 3485
rect 2665 3415 2685 3435
rect 2665 3365 2685 3385
rect 2665 3315 2685 3335
rect 2665 3265 2685 3285
rect 2665 3215 2685 3235
rect 2665 3165 2685 3185
rect 2665 3115 2685 3135
rect 1865 715 1885 735
rect 1865 665 1885 685
rect 1865 615 1885 635
rect 1865 565 1885 585
rect 1865 515 1885 535
rect 1865 465 1885 485
rect 1865 415 1885 435
rect 1865 365 1885 385
rect 1865 315 1885 335
rect 1865 265 1885 285
rect 1965 715 1985 735
rect 1965 665 1985 685
rect 1965 615 1985 635
rect 1965 565 1985 585
rect 1965 515 1985 535
rect 1965 465 1985 485
rect 1965 415 1985 435
rect 1965 365 1985 385
rect 1965 315 1985 335
rect 1965 265 1985 285
rect 2065 715 2085 735
rect 2065 665 2085 685
rect 2065 615 2085 635
rect 2065 565 2085 585
rect 2065 515 2085 535
rect 2065 465 2085 485
rect 2065 415 2085 435
rect 2065 365 2085 385
rect 2065 315 2085 335
rect 2065 265 2085 285
rect 2165 715 2185 735
rect 2165 665 2185 685
rect 2165 615 2185 635
rect 2165 565 2185 585
rect 2165 515 2185 535
rect 2165 465 2185 485
rect 2165 415 2185 435
rect 2165 365 2185 385
rect 2165 315 2185 335
rect 2165 265 2185 285
rect 2265 715 2285 735
rect 2265 665 2285 685
rect 2265 615 2285 635
rect 2265 565 2285 585
rect 2265 515 2285 535
rect 2265 465 2285 485
rect 2265 415 2285 435
rect 2265 365 2285 385
rect 2265 315 2285 335
rect 2265 265 2285 285
rect 2365 715 2385 735
rect 2365 665 2385 685
rect 2365 615 2385 635
rect 2365 565 2385 585
rect 2365 515 2385 535
rect 2365 465 2385 485
rect 2365 415 2385 435
rect 2365 365 2385 385
rect 2365 315 2385 335
rect 2365 265 2385 285
rect 2465 715 2485 735
rect 2465 665 2485 685
rect 2465 615 2485 635
rect 2465 565 2485 585
rect 2465 515 2485 535
rect 2465 465 2485 485
rect 2465 415 2485 435
rect 2465 365 2485 385
rect 2465 315 2485 335
rect 2465 265 2485 285
rect 2565 715 2585 735
rect 2565 665 2585 685
rect 2565 615 2585 635
rect 2565 565 2585 585
rect 2565 515 2585 535
rect 2565 465 2585 485
rect 2565 415 2585 435
rect 2565 365 2585 385
rect 2565 315 2585 335
rect 2565 265 2585 285
rect 2665 715 2685 735
rect 2665 665 2685 685
rect 2665 615 2685 635
rect 2665 565 2685 585
rect 2665 515 2685 535
rect 2665 465 2685 485
rect 2665 415 2685 435
rect 2665 365 2685 385
rect 2665 315 2685 335
rect 2665 265 2685 285
<< psubdiff >>
rect 1450 3835 3100 3850
rect 1450 3815 1465 3835
rect 1485 3815 1515 3835
rect 1535 3815 1565 3835
rect 1585 3815 1615 3835
rect 1635 3815 1665 3835
rect 1685 3815 1715 3835
rect 1735 3815 1765 3835
rect 1785 3815 1815 3835
rect 1835 3815 1865 3835
rect 1885 3815 1915 3835
rect 1935 3815 1965 3835
rect 1985 3815 2015 3835
rect 2035 3815 2065 3835
rect 2085 3815 2115 3835
rect 2135 3815 2165 3835
rect 2185 3815 2215 3835
rect 2235 3815 2265 3835
rect 2285 3815 2315 3835
rect 2335 3815 2365 3835
rect 2385 3815 2415 3835
rect 2435 3815 2465 3835
rect 2485 3815 2515 3835
rect 2535 3815 2565 3835
rect 2585 3815 2615 3835
rect 2635 3815 2665 3835
rect 2685 3815 2715 3835
rect 2735 3815 2765 3835
rect 2785 3815 2815 3835
rect 2835 3815 2865 3835
rect 2885 3815 2915 3835
rect 2935 3815 2965 3835
rect 2985 3815 3015 3835
rect 3035 3815 3065 3835
rect 3085 3815 3100 3835
rect 1450 3800 3100 3815
rect 1450 3785 1500 3800
rect 1450 3765 1465 3785
rect 1485 3765 1500 3785
rect 1450 3735 1500 3765
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1450 3685 1500 3715
rect 3050 3785 3100 3800
rect 3050 3765 3065 3785
rect 3085 3765 3100 3785
rect 3050 3735 3100 3765
rect 3050 3715 3065 3735
rect 3085 3715 3100 3735
rect 1450 3665 1465 3685
rect 1485 3665 1500 3685
rect 1450 3635 1500 3665
rect 1450 3615 1465 3635
rect 1485 3615 1500 3635
rect 1450 3585 1500 3615
rect 1450 3565 1465 3585
rect 1485 3565 1500 3585
rect 1450 3535 1500 3565
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3285 1500 3315
rect 1450 3265 1465 3285
rect 1485 3265 1500 3285
rect 1450 3235 1500 3265
rect 1450 3215 1465 3235
rect 1485 3215 1500 3235
rect 1450 3185 1500 3215
rect 1450 3165 1465 3185
rect 1485 3165 1500 3185
rect 1450 3135 1500 3165
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3085 1500 3115
rect 1450 3065 1465 3085
rect 1485 3065 1500 3085
rect 1450 3035 1500 3065
rect 1450 3015 1465 3035
rect 1485 3015 1500 3035
rect 1450 2985 1500 3015
rect 1450 2965 1465 2985
rect 1485 2965 1500 2985
rect 1450 2935 1500 2965
rect 1450 2915 1465 2935
rect 1485 2915 1500 2935
rect 1450 2885 1500 2915
rect 1450 2865 1465 2885
rect 1485 2865 1500 2885
rect 1450 2835 1500 2865
rect 1450 2815 1465 2835
rect 1485 2815 1500 2835
rect 1450 2785 1500 2815
rect 1450 2765 1465 2785
rect 1485 2765 1500 2785
rect 1450 2735 1500 2765
rect 1450 2715 1465 2735
rect 1485 2715 1500 2735
rect 1450 2685 1500 2715
rect 1450 2665 1465 2685
rect 1485 2665 1500 2685
rect 1450 2635 1500 2665
rect 1450 2615 1465 2635
rect 1485 2615 1500 2635
rect 1450 2585 1500 2615
rect 1450 2565 1465 2585
rect 1485 2565 1500 2585
rect 1450 2535 1500 2565
rect 1450 2515 1465 2535
rect 1485 2515 1500 2535
rect 1450 2485 1500 2515
rect 1450 2465 1465 2485
rect 1485 2465 1500 2485
rect 1450 2435 1500 2465
rect 1450 2415 1465 2435
rect 1485 2415 1500 2435
rect 1450 2385 1500 2415
rect 1450 2365 1465 2385
rect 1485 2365 1500 2385
rect 1450 2335 1500 2365
rect 1450 2315 1465 2335
rect 1485 2315 1500 2335
rect 1450 2285 1500 2315
rect 1450 2265 1465 2285
rect 1485 2265 1500 2285
rect 1450 2235 1500 2265
rect 1450 2215 1465 2235
rect 1485 2215 1500 2235
rect 1450 2185 1500 2215
rect 1450 2165 1465 2185
rect 1485 2165 1500 2185
rect 1450 2135 1500 2165
rect 1450 2115 1465 2135
rect 1485 2115 1500 2135
rect 1450 2085 1500 2115
rect 1450 2065 1465 2085
rect 1485 2065 1500 2085
rect 1450 2035 1500 2065
rect 1450 2015 1465 2035
rect 1485 2015 1500 2035
rect 1450 1985 1500 2015
rect 1450 1965 1465 1985
rect 1485 1965 1500 1985
rect 1450 1935 1500 1965
rect 1450 1915 1465 1935
rect 1485 1915 1500 1935
rect 1450 1885 1500 1915
rect 1450 1865 1465 1885
rect 1485 1865 1500 1885
rect 1450 1835 1500 1865
rect 1450 1815 1465 1835
rect 1485 1815 1500 1835
rect 1450 1785 1500 1815
rect 1450 1765 1465 1785
rect 1485 1765 1500 1785
rect 1450 1735 1500 1765
rect 1450 1715 1465 1735
rect 1485 1715 1500 1735
rect 1450 1685 1500 1715
rect 1450 1665 1465 1685
rect 1485 1665 1500 1685
rect 1450 1635 1500 1665
rect 1450 1615 1465 1635
rect 1485 1615 1500 1635
rect 1450 1585 1500 1615
rect 1450 1565 1465 1585
rect 1485 1565 1500 1585
rect 1450 1535 1500 1565
rect 1450 1515 1465 1535
rect 1485 1515 1500 1535
rect 1450 1485 1500 1515
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 935 1500 965
rect 1450 915 1465 935
rect 1485 915 1500 935
rect 1450 885 1500 915
rect 1450 865 1465 885
rect 1485 865 1500 885
rect 1450 835 1500 865
rect 1450 815 1465 835
rect 1485 815 1500 835
rect 1450 785 1500 815
rect 1450 765 1465 785
rect 1485 765 1500 785
rect 1450 735 1500 765
rect 1450 715 1465 735
rect 1485 715 1500 735
rect 1450 685 1500 715
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 135 1500 165
rect 1750 2785 2800 2800
rect 1750 2765 1765 2785
rect 1785 2765 1815 2785
rect 1835 2765 1865 2785
rect 1885 2765 1915 2785
rect 1935 2765 1965 2785
rect 1985 2765 2015 2785
rect 2035 2765 2065 2785
rect 2085 2765 2115 2785
rect 2135 2765 2165 2785
rect 2185 2765 2215 2785
rect 2235 2765 2265 2785
rect 2285 2765 2315 2785
rect 2335 2765 2365 2785
rect 2385 2765 2415 2785
rect 2435 2765 2465 2785
rect 2485 2765 2515 2785
rect 2535 2765 2565 2785
rect 2585 2765 2615 2785
rect 2635 2765 2665 2785
rect 2685 2765 2715 2785
rect 2735 2765 2765 2785
rect 2785 2765 2800 2785
rect 1750 2750 2800 2765
rect 1750 2735 1800 2750
rect 1750 2715 1765 2735
rect 1785 2715 1800 2735
rect 2750 2735 2800 2750
rect 2750 2715 2765 2735
rect 2785 2715 2800 2735
rect 1750 2685 1800 2715
rect 1750 2665 1765 2685
rect 1785 2665 1800 2685
rect 1750 2635 1800 2665
rect 1750 2615 1765 2635
rect 1785 2615 1800 2635
rect 1750 2585 1800 2615
rect 1750 2565 1765 2585
rect 1785 2565 1800 2585
rect 1750 2535 1800 2565
rect 1750 2515 1765 2535
rect 1785 2515 1800 2535
rect 1750 2485 1800 2515
rect 1750 2465 1765 2485
rect 1785 2465 1800 2485
rect 1750 2435 1800 2465
rect 1750 2415 1765 2435
rect 1785 2415 1800 2435
rect 1750 2385 1800 2415
rect 1750 2365 1765 2385
rect 1785 2365 1800 2385
rect 1750 2335 1800 2365
rect 1750 2315 1765 2335
rect 1785 2315 1800 2335
rect 1750 2285 1800 2315
rect 1750 2265 1765 2285
rect 1785 2265 1800 2285
rect 1750 2235 1800 2265
rect 1750 2215 1765 2235
rect 1785 2215 1800 2235
rect 1750 2185 1800 2215
rect 1750 2165 1765 2185
rect 1785 2165 1800 2185
rect 1750 2135 1800 2165
rect 1750 2115 1765 2135
rect 1785 2115 1800 2135
rect 1750 2085 1800 2115
rect 1750 2065 1765 2085
rect 1785 2065 1800 2085
rect 1750 2035 1800 2065
rect 1750 2015 1765 2035
rect 1785 2015 1800 2035
rect 1750 1985 1800 2015
rect 2750 2685 2800 2715
rect 2750 2665 2765 2685
rect 2785 2665 2800 2685
rect 2750 2635 2800 2665
rect 2750 2615 2765 2635
rect 2785 2615 2800 2635
rect 2750 2585 2800 2615
rect 2750 2565 2765 2585
rect 2785 2565 2800 2585
rect 2750 2535 2800 2565
rect 2750 2515 2765 2535
rect 2785 2515 2800 2535
rect 2750 2485 2800 2515
rect 2750 2465 2765 2485
rect 2785 2465 2800 2485
rect 2750 2435 2800 2465
rect 2750 2415 2765 2435
rect 2785 2415 2800 2435
rect 2750 2385 2800 2415
rect 2750 2365 2765 2385
rect 2785 2365 2800 2385
rect 2750 2335 2800 2365
rect 2750 2315 2765 2335
rect 2785 2315 2800 2335
rect 2750 2285 2800 2315
rect 2750 2265 2765 2285
rect 2785 2265 2800 2285
rect 2750 2235 2800 2265
rect 2750 2215 2765 2235
rect 2785 2215 2800 2235
rect 2750 2185 2800 2215
rect 2750 2165 2765 2185
rect 2785 2165 2800 2185
rect 2750 2135 2800 2165
rect 2750 2115 2765 2135
rect 2785 2115 2800 2135
rect 2750 2085 2800 2115
rect 2750 2065 2765 2085
rect 2785 2065 2800 2085
rect 2750 2035 2800 2065
rect 2750 2015 2765 2035
rect 2785 2015 2800 2035
rect 1750 1965 1765 1985
rect 1785 1965 1800 1985
rect 1750 1935 1800 1965
rect 1750 1915 1765 1935
rect 1785 1915 1800 1935
rect 1750 1885 1800 1915
rect 1750 1865 1765 1885
rect 1785 1865 1800 1885
rect 1750 1835 1800 1865
rect 2750 1985 2800 2015
rect 2750 1965 2765 1985
rect 2785 1965 2800 1985
rect 2750 1935 2800 1965
rect 2750 1915 2765 1935
rect 2785 1915 2800 1935
rect 2750 1885 2800 1915
rect 2750 1865 2765 1885
rect 2785 1865 2800 1885
rect 1750 1815 1765 1835
rect 1785 1815 1800 1835
rect 1750 1785 1800 1815
rect 1750 1765 1765 1785
rect 1785 1765 1800 1785
rect 1750 1735 1800 1765
rect 1750 1715 1765 1735
rect 1785 1715 1800 1735
rect 1750 1685 1800 1715
rect 1750 1665 1765 1685
rect 1785 1665 1800 1685
rect 1750 1635 1800 1665
rect 1750 1615 1765 1635
rect 1785 1615 1800 1635
rect 1750 1585 1800 1615
rect 1750 1565 1765 1585
rect 1785 1565 1800 1585
rect 1750 1535 1800 1565
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1750 1485 1800 1515
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 2750 1835 2800 1865
rect 2750 1815 2765 1835
rect 2785 1815 2800 1835
rect 2750 1785 2800 1815
rect 2750 1765 2765 1785
rect 2785 1765 2800 1785
rect 2750 1735 2800 1765
rect 2750 1715 2765 1735
rect 2785 1715 2800 1735
rect 2750 1685 2800 1715
rect 2750 1665 2765 1685
rect 2785 1665 2800 1685
rect 2750 1635 2800 1665
rect 2750 1615 2765 1635
rect 2785 1615 2800 1635
rect 2750 1585 2800 1615
rect 2750 1565 2765 1585
rect 2785 1565 2800 1585
rect 2750 1535 2800 1565
rect 2750 1515 2765 1535
rect 2785 1515 2800 1535
rect 2750 1485 2800 1515
rect 2750 1465 2765 1485
rect 2785 1465 2800 1485
rect 2750 1435 2800 1465
rect 2750 1415 2765 1435
rect 2785 1415 2800 1435
rect 2750 1385 2800 1415
rect 2750 1365 2765 1385
rect 2785 1365 2800 1385
rect 2750 1335 2800 1365
rect 2750 1315 2765 1335
rect 2785 1315 2800 1335
rect 2750 1285 2800 1315
rect 2750 1265 2765 1285
rect 2785 1265 2800 1285
rect 2750 1235 2800 1265
rect 2750 1215 2765 1235
rect 2785 1215 2800 1235
rect 2750 1185 2800 1215
rect 2750 1165 2765 1185
rect 2785 1165 2800 1185
rect 2750 1135 2800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1100 1800 1115
rect 2750 1115 2765 1135
rect 2785 1115 2800 1135
rect 2750 1100 2800 1115
rect 1750 1085 2800 1100
rect 1750 1065 1765 1085
rect 1785 1065 1815 1085
rect 1835 1065 1865 1085
rect 1885 1065 1915 1085
rect 1935 1065 1965 1085
rect 1985 1065 2015 1085
rect 2035 1065 2065 1085
rect 2085 1065 2115 1085
rect 2135 1065 2165 1085
rect 2185 1065 2215 1085
rect 2235 1065 2265 1085
rect 2285 1065 2315 1085
rect 2335 1065 2365 1085
rect 2385 1065 2415 1085
rect 2435 1065 2465 1085
rect 2485 1065 2515 1085
rect 2535 1065 2565 1085
rect 2585 1065 2615 1085
rect 2635 1065 2665 1085
rect 2685 1065 2715 1085
rect 2735 1065 2765 1085
rect 2785 1065 2800 1085
rect 1750 1050 2800 1065
rect 3050 3685 3100 3715
rect 3050 3665 3065 3685
rect 3085 3665 3100 3685
rect 3050 3635 3100 3665
rect 3050 3615 3065 3635
rect 3085 3615 3100 3635
rect 3050 3585 3100 3615
rect 3050 3565 3065 3585
rect 3085 3565 3100 3585
rect 3050 3535 3100 3565
rect 3050 3515 3065 3535
rect 3085 3515 3100 3535
rect 3050 3485 3100 3515
rect 3050 3465 3065 3485
rect 3085 3465 3100 3485
rect 3050 3435 3100 3465
rect 3050 3415 3065 3435
rect 3085 3415 3100 3435
rect 3050 3385 3100 3415
rect 3050 3365 3065 3385
rect 3085 3365 3100 3385
rect 3050 3335 3100 3365
rect 3050 3315 3065 3335
rect 3085 3315 3100 3335
rect 3050 3285 3100 3315
rect 3050 3265 3065 3285
rect 3085 3265 3100 3285
rect 3050 3235 3100 3265
rect 3050 3215 3065 3235
rect 3085 3215 3100 3235
rect 3050 3185 3100 3215
rect 3050 3165 3065 3185
rect 3085 3165 3100 3185
rect 3050 3135 3100 3165
rect 3050 3115 3065 3135
rect 3085 3115 3100 3135
rect 3050 3085 3100 3115
rect 3050 3065 3065 3085
rect 3085 3065 3100 3085
rect 3050 3035 3100 3065
rect 3050 3015 3065 3035
rect 3085 3015 3100 3035
rect 3050 2985 3100 3015
rect 3050 2965 3065 2985
rect 3085 2965 3100 2985
rect 3050 2935 3100 2965
rect 3050 2915 3065 2935
rect 3085 2915 3100 2935
rect 3050 2885 3100 2915
rect 3050 2865 3065 2885
rect 3085 2865 3100 2885
rect 3050 2835 3100 2865
rect 3050 2815 3065 2835
rect 3085 2815 3100 2835
rect 3050 2785 3100 2815
rect 3050 2765 3065 2785
rect 3085 2765 3100 2785
rect 3050 2735 3100 2765
rect 3050 2715 3065 2735
rect 3085 2715 3100 2735
rect 3050 2685 3100 2715
rect 3050 2665 3065 2685
rect 3085 2665 3100 2685
rect 3050 2635 3100 2665
rect 3050 2615 3065 2635
rect 3085 2615 3100 2635
rect 3050 2585 3100 2615
rect 3050 2565 3065 2585
rect 3085 2565 3100 2585
rect 3050 2535 3100 2565
rect 3050 2515 3065 2535
rect 3085 2515 3100 2535
rect 3050 2485 3100 2515
rect 3050 2465 3065 2485
rect 3085 2465 3100 2485
rect 3050 2435 3100 2465
rect 3050 2415 3065 2435
rect 3085 2415 3100 2435
rect 3050 2385 3100 2415
rect 3050 2365 3065 2385
rect 3085 2365 3100 2385
rect 3050 2335 3100 2365
rect 3050 2315 3065 2335
rect 3085 2315 3100 2335
rect 3050 2285 3100 2315
rect 3050 2265 3065 2285
rect 3085 2265 3100 2285
rect 3050 2235 3100 2265
rect 3050 2215 3065 2235
rect 3085 2215 3100 2235
rect 3050 2185 3100 2215
rect 3050 2165 3065 2185
rect 3085 2165 3100 2185
rect 3050 2135 3100 2165
rect 3050 2115 3065 2135
rect 3085 2115 3100 2135
rect 3050 2085 3100 2115
rect 3050 2065 3065 2085
rect 3085 2065 3100 2085
rect 3050 2035 3100 2065
rect 3050 2015 3065 2035
rect 3085 2015 3100 2035
rect 3050 1985 3100 2015
rect 3050 1965 3065 1985
rect 3085 1965 3100 1985
rect 3050 1935 3100 1965
rect 3050 1915 3065 1935
rect 3085 1915 3100 1935
rect 3050 1885 3100 1915
rect 3050 1865 3065 1885
rect 3085 1865 3100 1885
rect 3050 1835 3100 1865
rect 3050 1815 3065 1835
rect 3085 1815 3100 1835
rect 3050 1785 3100 1815
rect 3050 1765 3065 1785
rect 3085 1765 3100 1785
rect 3050 1735 3100 1765
rect 3050 1715 3065 1735
rect 3085 1715 3100 1735
rect 3050 1685 3100 1715
rect 3050 1665 3065 1685
rect 3085 1665 3100 1685
rect 3050 1635 3100 1665
rect 3050 1615 3065 1635
rect 3085 1615 3100 1635
rect 3050 1585 3100 1615
rect 3050 1565 3065 1585
rect 3085 1565 3100 1585
rect 3050 1535 3100 1565
rect 3050 1515 3065 1535
rect 3085 1515 3100 1535
rect 3050 1485 3100 1515
rect 3050 1465 3065 1485
rect 3085 1465 3100 1485
rect 3050 1435 3100 1465
rect 3050 1415 3065 1435
rect 3085 1415 3100 1435
rect 3050 1385 3100 1415
rect 3050 1365 3065 1385
rect 3085 1365 3100 1385
rect 3050 1335 3100 1365
rect 3050 1315 3065 1335
rect 3085 1315 3100 1335
rect 3050 1285 3100 1315
rect 3050 1265 3065 1285
rect 3085 1265 3100 1285
rect 3050 1235 3100 1265
rect 3050 1215 3065 1235
rect 3085 1215 3100 1235
rect 3050 1185 3100 1215
rect 3050 1165 3065 1185
rect 3085 1165 3100 1185
rect 3050 1135 3100 1165
rect 3050 1115 3065 1135
rect 3085 1115 3100 1135
rect 3050 1085 3100 1115
rect 3050 1065 3065 1085
rect 3085 1065 3100 1085
rect 3050 1035 3100 1065
rect 3050 1015 3065 1035
rect 3085 1015 3100 1035
rect 3050 985 3100 1015
rect 3050 965 3065 985
rect 3085 965 3100 985
rect 3050 935 3100 965
rect 3050 915 3065 935
rect 3085 915 3100 935
rect 3050 885 3100 915
rect 3050 865 3065 885
rect 3085 865 3100 885
rect 3050 835 3100 865
rect 3050 815 3065 835
rect 3085 815 3100 835
rect 3050 785 3100 815
rect 3050 765 3065 785
rect 3085 765 3100 785
rect 3050 735 3100 765
rect 3050 715 3065 735
rect 3085 715 3100 735
rect 3050 685 3100 715
rect 3050 665 3065 685
rect 3085 665 3100 685
rect 3050 635 3100 665
rect 3050 615 3065 635
rect 3085 615 3100 635
rect 3050 585 3100 615
rect 3050 565 3065 585
rect 3085 565 3100 585
rect 3050 535 3100 565
rect 3050 515 3065 535
rect 3085 515 3100 535
rect 3050 485 3100 515
rect 3050 465 3065 485
rect 3085 465 3100 485
rect 3050 435 3100 465
rect 3050 415 3065 435
rect 3085 415 3100 435
rect 3050 385 3100 415
rect 3050 365 3065 385
rect 3085 365 3100 385
rect 3050 335 3100 365
rect 3050 315 3065 335
rect 3085 315 3100 335
rect 3050 285 3100 315
rect 3050 265 3065 285
rect 3085 265 3100 285
rect 3050 235 3100 265
rect 3050 215 3065 235
rect 3085 215 3100 235
rect 3050 185 3100 215
rect 3050 165 3065 185
rect 3085 165 3100 185
rect 1450 115 1465 135
rect 1485 115 1500 135
rect 1450 85 1500 115
rect 1450 65 1465 85
rect 1485 65 1500 85
rect 1450 50 1500 65
rect 3050 135 3100 165
rect 3050 115 3065 135
rect 3085 115 3100 135
rect 3050 85 3100 115
rect 3050 65 3065 85
rect 3085 65 3100 85
rect 3050 50 3100 65
rect 1450 35 3100 50
rect 1450 15 1465 35
rect 1485 15 1515 35
rect 1535 15 1565 35
rect 1585 15 1615 35
rect 1635 15 1665 35
rect 1685 15 1715 35
rect 1735 15 1765 35
rect 1785 15 1815 35
rect 1835 15 1865 35
rect 1885 15 1915 35
rect 1935 15 1965 35
rect 1985 15 2015 35
rect 2035 15 2065 35
rect 2085 15 2115 35
rect 2135 15 2165 35
rect 2185 15 2215 35
rect 2235 15 2265 35
rect 2285 15 2315 35
rect 2335 15 2365 35
rect 2385 15 2415 35
rect 2435 15 2465 35
rect 2485 15 2515 35
rect 2535 15 2565 35
rect 2585 15 2615 35
rect 2635 15 2665 35
rect 2685 15 2715 35
rect 2735 15 2765 35
rect 2785 15 2815 35
rect 2835 15 2865 35
rect 2885 15 2915 35
rect 2935 15 2965 35
rect 2985 15 3015 35
rect 3035 15 3065 35
rect 3085 15 3100 35
rect 1450 0 3100 15
<< nsubdiff >>
rect 1600 3685 2950 3700
rect 1600 3665 1615 3685
rect 1635 3665 1665 3685
rect 1685 3665 1715 3685
rect 1735 3665 1765 3685
rect 1785 3665 1815 3685
rect 1835 3665 1865 3685
rect 1885 3665 1915 3685
rect 1935 3665 1965 3685
rect 1985 3665 2015 3685
rect 2035 3665 2065 3685
rect 2085 3665 2115 3685
rect 2135 3665 2165 3685
rect 2185 3665 2215 3685
rect 2235 3665 2265 3685
rect 2285 3665 2315 3685
rect 2335 3665 2365 3685
rect 2385 3665 2415 3685
rect 2435 3665 2465 3685
rect 2485 3665 2515 3685
rect 2535 3665 2565 3685
rect 2585 3665 2615 3685
rect 2635 3665 2665 3685
rect 2685 3665 2715 3685
rect 2735 3665 2765 3685
rect 2785 3665 2815 3685
rect 2835 3665 2865 3685
rect 2885 3665 2915 3685
rect 2935 3665 2950 3685
rect 1600 3650 2950 3665
rect 1600 3635 1650 3650
rect 1600 3615 1615 3635
rect 1635 3615 1650 3635
rect 2900 3635 2950 3650
rect 2900 3615 2915 3635
rect 2935 3615 2950 3635
rect 1600 3585 1650 3615
rect 1600 3565 1615 3585
rect 1635 3565 1650 3585
rect 1600 3535 1650 3565
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3285 1650 3315
rect 1600 3265 1615 3285
rect 1635 3265 1650 3285
rect 1600 3235 1650 3265
rect 1600 3215 1615 3235
rect 1635 3215 1650 3235
rect 1600 3185 1650 3215
rect 1600 3165 1615 3185
rect 1635 3165 1650 3185
rect 1600 3135 1650 3165
rect 1600 3115 1615 3135
rect 1635 3115 1650 3135
rect 1600 3085 1650 3115
rect 2900 3585 2950 3615
rect 2900 3565 2915 3585
rect 2935 3565 2950 3585
rect 2900 3535 2950 3565
rect 2900 3515 2915 3535
rect 2935 3515 2950 3535
rect 2900 3485 2950 3515
rect 2900 3465 2915 3485
rect 2935 3465 2950 3485
rect 2900 3435 2950 3465
rect 2900 3415 2915 3435
rect 2935 3415 2950 3435
rect 2900 3385 2950 3415
rect 2900 3365 2915 3385
rect 2935 3365 2950 3385
rect 2900 3335 2950 3365
rect 2900 3315 2915 3335
rect 2935 3315 2950 3335
rect 2900 3285 2950 3315
rect 2900 3265 2915 3285
rect 2935 3265 2950 3285
rect 2900 3235 2950 3265
rect 2900 3215 2915 3235
rect 2935 3215 2950 3235
rect 2900 3185 2950 3215
rect 2900 3165 2915 3185
rect 2935 3165 2950 3185
rect 2900 3135 2950 3165
rect 2900 3115 2915 3135
rect 2935 3115 2950 3135
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1600 3035 1650 3065
rect 1600 3015 1615 3035
rect 1635 3015 1650 3035
rect 1600 2985 1650 3015
rect 2900 3085 2950 3115
rect 2900 3065 2915 3085
rect 2935 3065 2950 3085
rect 2900 3035 2950 3065
rect 2900 3015 2915 3035
rect 2935 3015 2950 3035
rect 1600 2965 1615 2985
rect 1635 2965 1650 2985
rect 1600 2950 1650 2965
rect 2900 2985 2950 3015
rect 2900 2965 2915 2985
rect 2935 2965 2950 2985
rect 2900 2950 2950 2965
rect 1600 2935 2950 2950
rect 1600 2915 1615 2935
rect 1635 2915 1665 2935
rect 1685 2915 1715 2935
rect 1735 2915 1765 2935
rect 1785 2915 1815 2935
rect 1835 2915 1865 2935
rect 1885 2915 1915 2935
rect 1935 2915 1965 2935
rect 1985 2915 2015 2935
rect 2035 2915 2065 2935
rect 2085 2915 2115 2935
rect 2135 2915 2165 2935
rect 2185 2915 2215 2935
rect 2235 2915 2265 2935
rect 2285 2915 2315 2935
rect 2335 2915 2365 2935
rect 2385 2915 2415 2935
rect 2435 2915 2465 2935
rect 2485 2915 2515 2935
rect 2535 2915 2565 2935
rect 2585 2915 2615 2935
rect 2635 2915 2665 2935
rect 2685 2915 2715 2935
rect 2735 2915 2765 2935
rect 2785 2915 2815 2935
rect 2835 2915 2865 2935
rect 2885 2915 2915 2935
rect 2935 2915 2950 2935
rect 1600 2900 2950 2915
rect 1600 2885 1650 2900
rect 1600 2865 1615 2885
rect 1635 2865 1650 2885
rect 1600 2835 1650 2865
rect 1600 2815 1615 2835
rect 1635 2815 1650 2835
rect 1600 2785 1650 2815
rect 2900 2885 2950 2900
rect 2900 2865 2915 2885
rect 2935 2865 2950 2885
rect 2900 2835 2950 2865
rect 2900 2815 2915 2835
rect 2935 2815 2950 2835
rect 1600 2765 1615 2785
rect 1635 2765 1650 2785
rect 1600 2735 1650 2765
rect 1600 2715 1615 2735
rect 1635 2715 1650 2735
rect 1600 2685 1650 2715
rect 1600 2665 1615 2685
rect 1635 2665 1650 2685
rect 1600 2635 1650 2665
rect 1600 2615 1615 2635
rect 1635 2615 1650 2635
rect 1600 2585 1650 2615
rect 1600 2565 1615 2585
rect 1635 2565 1650 2585
rect 1600 2535 1650 2565
rect 1600 2515 1615 2535
rect 1635 2515 1650 2535
rect 1600 2485 1650 2515
rect 1600 2465 1615 2485
rect 1635 2465 1650 2485
rect 1600 2435 1650 2465
rect 1600 2415 1615 2435
rect 1635 2415 1650 2435
rect 1600 2385 1650 2415
rect 1600 2365 1615 2385
rect 1635 2365 1650 2385
rect 1600 2335 1650 2365
rect 1600 2315 1615 2335
rect 1635 2315 1650 2335
rect 1600 2285 1650 2315
rect 1600 2265 1615 2285
rect 1635 2265 1650 2285
rect 1600 2235 1650 2265
rect 1600 2215 1615 2235
rect 1635 2215 1650 2235
rect 1600 2185 1650 2215
rect 1600 2165 1615 2185
rect 1635 2165 1650 2185
rect 1600 2135 1650 2165
rect 1600 2115 1615 2135
rect 1635 2115 1650 2135
rect 1600 2085 1650 2115
rect 1600 2065 1615 2085
rect 1635 2065 1650 2085
rect 1600 2035 1650 2065
rect 1600 2015 1615 2035
rect 1635 2015 1650 2035
rect 1600 1985 1650 2015
rect 1600 1965 1615 1985
rect 1635 1965 1650 1985
rect 1600 1935 1650 1965
rect 1600 1915 1615 1935
rect 1635 1915 1650 1935
rect 1600 1885 1650 1915
rect 1600 1865 1615 1885
rect 1635 1865 1650 1885
rect 1600 1835 1650 1865
rect 1600 1815 1615 1835
rect 1635 1815 1650 1835
rect 1600 1785 1650 1815
rect 1600 1765 1615 1785
rect 1635 1765 1650 1785
rect 1600 1735 1650 1765
rect 1600 1715 1615 1735
rect 1635 1715 1650 1735
rect 1600 1685 1650 1715
rect 1600 1665 1615 1685
rect 1635 1665 1650 1685
rect 1600 1635 1650 1665
rect 1600 1615 1615 1635
rect 1635 1615 1650 1635
rect 1600 1585 1650 1615
rect 1600 1565 1615 1585
rect 1635 1565 1650 1585
rect 1600 1535 1650 1565
rect 1600 1515 1615 1535
rect 1635 1515 1650 1535
rect 1600 1485 1650 1515
rect 1600 1465 1615 1485
rect 1635 1465 1650 1485
rect 1600 1435 1650 1465
rect 1600 1415 1615 1435
rect 1635 1415 1650 1435
rect 1600 1385 1650 1415
rect 1600 1365 1615 1385
rect 1635 1365 1650 1385
rect 1600 1335 1650 1365
rect 1600 1315 1615 1335
rect 1635 1315 1650 1335
rect 1600 1285 1650 1315
rect 1600 1265 1615 1285
rect 1635 1265 1650 1285
rect 1600 1235 1650 1265
rect 1600 1215 1615 1235
rect 1635 1215 1650 1235
rect 1600 1185 1650 1215
rect 1600 1165 1615 1185
rect 1635 1165 1650 1185
rect 1600 1135 1650 1165
rect 1600 1115 1615 1135
rect 1635 1115 1650 1135
rect 1600 1085 1650 1115
rect 1600 1065 1615 1085
rect 1635 1065 1650 1085
rect 1600 1035 1650 1065
rect 2900 2785 2950 2815
rect 2900 2765 2915 2785
rect 2935 2765 2950 2785
rect 2900 2735 2950 2765
rect 2900 2715 2915 2735
rect 2935 2715 2950 2735
rect 2900 2685 2950 2715
rect 2900 2665 2915 2685
rect 2935 2665 2950 2685
rect 2900 2635 2950 2665
rect 2900 2615 2915 2635
rect 2935 2615 2950 2635
rect 2900 2585 2950 2615
rect 2900 2565 2915 2585
rect 2935 2565 2950 2585
rect 2900 2535 2950 2565
rect 2900 2515 2915 2535
rect 2935 2515 2950 2535
rect 2900 2485 2950 2515
rect 2900 2465 2915 2485
rect 2935 2465 2950 2485
rect 2900 2435 2950 2465
rect 2900 2415 2915 2435
rect 2935 2415 2950 2435
rect 2900 2385 2950 2415
rect 2900 2365 2915 2385
rect 2935 2365 2950 2385
rect 2900 2335 2950 2365
rect 2900 2315 2915 2335
rect 2935 2315 2950 2335
rect 2900 2285 2950 2315
rect 2900 2265 2915 2285
rect 2935 2265 2950 2285
rect 2900 2235 2950 2265
rect 2900 2215 2915 2235
rect 2935 2215 2950 2235
rect 2900 2185 2950 2215
rect 2900 2165 2915 2185
rect 2935 2165 2950 2185
rect 2900 2135 2950 2165
rect 2900 2115 2915 2135
rect 2935 2115 2950 2135
rect 2900 2085 2950 2115
rect 2900 2065 2915 2085
rect 2935 2065 2950 2085
rect 2900 2035 2950 2065
rect 2900 2015 2915 2035
rect 2935 2015 2950 2035
rect 2900 1985 2950 2015
rect 2900 1965 2915 1985
rect 2935 1965 2950 1985
rect 2900 1935 2950 1965
rect 2900 1915 2915 1935
rect 2935 1915 2950 1935
rect 2900 1885 2950 1915
rect 2900 1865 2915 1885
rect 2935 1865 2950 1885
rect 2900 1835 2950 1865
rect 2900 1815 2915 1835
rect 2935 1815 2950 1835
rect 2900 1785 2950 1815
rect 2900 1765 2915 1785
rect 2935 1765 2950 1785
rect 2900 1735 2950 1765
rect 2900 1715 2915 1735
rect 2935 1715 2950 1735
rect 2900 1685 2950 1715
rect 2900 1665 2915 1685
rect 2935 1665 2950 1685
rect 2900 1635 2950 1665
rect 2900 1615 2915 1635
rect 2935 1615 2950 1635
rect 2900 1585 2950 1615
rect 2900 1565 2915 1585
rect 2935 1565 2950 1585
rect 2900 1535 2950 1565
rect 2900 1515 2915 1535
rect 2935 1515 2950 1535
rect 2900 1485 2950 1515
rect 2900 1465 2915 1485
rect 2935 1465 2950 1485
rect 2900 1435 2950 1465
rect 2900 1415 2915 1435
rect 2935 1415 2950 1435
rect 2900 1385 2950 1415
rect 2900 1365 2915 1385
rect 2935 1365 2950 1385
rect 2900 1335 2950 1365
rect 2900 1315 2915 1335
rect 2935 1315 2950 1335
rect 2900 1285 2950 1315
rect 2900 1265 2915 1285
rect 2935 1265 2950 1285
rect 2900 1235 2950 1265
rect 2900 1215 2915 1235
rect 2935 1215 2950 1235
rect 2900 1185 2950 1215
rect 2900 1165 2915 1185
rect 2935 1165 2950 1185
rect 2900 1135 2950 1165
rect 2900 1115 2915 1135
rect 2935 1115 2950 1135
rect 2900 1085 2950 1115
rect 2900 1065 2915 1085
rect 2935 1065 2950 1085
rect 1600 1015 1615 1035
rect 1635 1015 1650 1035
rect 1600 985 1650 1015
rect 1600 965 1615 985
rect 1635 965 1650 985
rect 1600 950 1650 965
rect 2900 1035 2950 1065
rect 2900 1015 2915 1035
rect 2935 1015 2950 1035
rect 2900 985 2950 1015
rect 2900 965 2915 985
rect 2935 965 2950 985
rect 2900 950 2950 965
rect 1600 935 2950 950
rect 1600 915 1615 935
rect 1635 915 1665 935
rect 1685 915 1715 935
rect 1735 915 1765 935
rect 1785 915 1815 935
rect 1835 915 1865 935
rect 1885 915 1915 935
rect 1935 915 1965 935
rect 1985 915 2015 935
rect 2035 915 2065 935
rect 2085 915 2115 935
rect 2135 915 2165 935
rect 2185 915 2215 935
rect 2235 915 2265 935
rect 2285 915 2315 935
rect 2335 915 2365 935
rect 2385 915 2415 935
rect 2435 915 2465 935
rect 2485 915 2515 935
rect 2535 915 2565 935
rect 2585 915 2615 935
rect 2635 915 2665 935
rect 2685 915 2715 935
rect 2735 915 2765 935
rect 2785 915 2815 935
rect 2835 915 2865 935
rect 2885 915 2915 935
rect 2935 915 2950 935
rect 1600 900 2950 915
rect 1600 885 1650 900
rect 1600 865 1615 885
rect 1635 865 1650 885
rect 1600 835 1650 865
rect 2900 885 2950 900
rect 2900 865 2915 885
rect 2935 865 2950 885
rect 1600 815 1615 835
rect 1635 815 1650 835
rect 1600 785 1650 815
rect 1600 765 1615 785
rect 1635 765 1650 785
rect 1600 735 1650 765
rect 2900 835 2950 865
rect 2900 815 2915 835
rect 2935 815 2950 835
rect 2900 785 2950 815
rect 2900 765 2915 785
rect 2935 765 2950 785
rect 1600 715 1615 735
rect 1635 715 1650 735
rect 1600 685 1650 715
rect 1600 665 1615 685
rect 1635 665 1650 685
rect 1600 635 1650 665
rect 1600 615 1615 635
rect 1635 615 1650 635
rect 1600 585 1650 615
rect 1600 565 1615 585
rect 1635 565 1650 585
rect 1600 535 1650 565
rect 1600 515 1615 535
rect 1635 515 1650 535
rect 1600 485 1650 515
rect 1600 465 1615 485
rect 1635 465 1650 485
rect 1600 435 1650 465
rect 1600 415 1615 435
rect 1635 415 1650 435
rect 1600 385 1650 415
rect 1600 365 1615 385
rect 1635 365 1650 385
rect 1600 335 1650 365
rect 1600 315 1615 335
rect 1635 315 1650 335
rect 1600 285 1650 315
rect 1600 265 1615 285
rect 1635 265 1650 285
rect 1600 235 1650 265
rect 2900 735 2950 765
rect 2900 715 2915 735
rect 2935 715 2950 735
rect 2900 685 2950 715
rect 2900 665 2915 685
rect 2935 665 2950 685
rect 2900 635 2950 665
rect 2900 615 2915 635
rect 2935 615 2950 635
rect 2900 585 2950 615
rect 2900 565 2915 585
rect 2935 565 2950 585
rect 2900 535 2950 565
rect 2900 515 2915 535
rect 2935 515 2950 535
rect 2900 485 2950 515
rect 2900 465 2915 485
rect 2935 465 2950 485
rect 2900 435 2950 465
rect 2900 415 2915 435
rect 2935 415 2950 435
rect 2900 385 2950 415
rect 2900 365 2915 385
rect 2935 365 2950 385
rect 2900 335 2950 365
rect 2900 315 2915 335
rect 2935 315 2950 335
rect 2900 285 2950 315
rect 2900 265 2915 285
rect 2935 265 2950 285
rect 2900 235 2950 265
rect 1600 215 1615 235
rect 1635 215 1650 235
rect 1600 200 1650 215
rect 2900 215 2915 235
rect 2935 215 2950 235
rect 2900 200 2950 215
rect 1600 185 2950 200
rect 1600 165 1615 185
rect 1635 165 1665 185
rect 1685 165 1715 185
rect 1735 165 1765 185
rect 1785 165 1815 185
rect 1835 165 1865 185
rect 1885 165 1915 185
rect 1935 165 1965 185
rect 1985 165 2015 185
rect 2035 165 2065 185
rect 2085 165 2115 185
rect 2135 165 2165 185
rect 2185 165 2215 185
rect 2235 165 2265 185
rect 2285 165 2315 185
rect 2335 165 2365 185
rect 2385 165 2415 185
rect 2435 165 2465 185
rect 2485 165 2515 185
rect 2535 165 2565 185
rect 2585 165 2615 185
rect 2635 165 2665 185
rect 2685 165 2715 185
rect 2735 165 2765 185
rect 2785 165 2815 185
rect 2835 165 2865 185
rect 2885 165 2915 185
rect 2935 165 2950 185
rect 1600 150 2950 165
<< psubdiffcont >>
rect 1465 3815 1485 3835
rect 1515 3815 1535 3835
rect 1565 3815 1585 3835
rect 1615 3815 1635 3835
rect 1665 3815 1685 3835
rect 1715 3815 1735 3835
rect 1765 3815 1785 3835
rect 1815 3815 1835 3835
rect 1865 3815 1885 3835
rect 1915 3815 1935 3835
rect 1965 3815 1985 3835
rect 2015 3815 2035 3835
rect 2065 3815 2085 3835
rect 2115 3815 2135 3835
rect 2165 3815 2185 3835
rect 2215 3815 2235 3835
rect 2265 3815 2285 3835
rect 2315 3815 2335 3835
rect 2365 3815 2385 3835
rect 2415 3815 2435 3835
rect 2465 3815 2485 3835
rect 2515 3815 2535 3835
rect 2565 3815 2585 3835
rect 2615 3815 2635 3835
rect 2665 3815 2685 3835
rect 2715 3815 2735 3835
rect 2765 3815 2785 3835
rect 2815 3815 2835 3835
rect 2865 3815 2885 3835
rect 2915 3815 2935 3835
rect 2965 3815 2985 3835
rect 3015 3815 3035 3835
rect 3065 3815 3085 3835
rect 1465 3765 1485 3785
rect 1465 3715 1485 3735
rect 3065 3765 3085 3785
rect 3065 3715 3085 3735
rect 1465 3665 1485 3685
rect 1465 3615 1485 3635
rect 1465 3565 1485 3585
rect 1465 3515 1485 3535
rect 1465 3465 1485 3485
rect 1465 3415 1485 3435
rect 1465 3365 1485 3385
rect 1465 3315 1485 3335
rect 1465 3265 1485 3285
rect 1465 3215 1485 3235
rect 1465 3165 1485 3185
rect 1465 3115 1485 3135
rect 1465 3065 1485 3085
rect 1465 3015 1485 3035
rect 1465 2965 1485 2985
rect 1465 2915 1485 2935
rect 1465 2865 1485 2885
rect 1465 2815 1485 2835
rect 1465 2765 1485 2785
rect 1465 2715 1485 2735
rect 1465 2665 1485 2685
rect 1465 2615 1485 2635
rect 1465 2565 1485 2585
rect 1465 2515 1485 2535
rect 1465 2465 1485 2485
rect 1465 2415 1485 2435
rect 1465 2365 1485 2385
rect 1465 2315 1485 2335
rect 1465 2265 1485 2285
rect 1465 2215 1485 2235
rect 1465 2165 1485 2185
rect 1465 2115 1485 2135
rect 1465 2065 1485 2085
rect 1465 2015 1485 2035
rect 1465 1965 1485 1985
rect 1465 1915 1485 1935
rect 1465 1865 1485 1885
rect 1465 1815 1485 1835
rect 1465 1765 1485 1785
rect 1465 1715 1485 1735
rect 1465 1665 1485 1685
rect 1465 1615 1485 1635
rect 1465 1565 1485 1585
rect 1465 1515 1485 1535
rect 1465 1465 1485 1485
rect 1465 1415 1485 1435
rect 1465 1365 1485 1385
rect 1465 1315 1485 1335
rect 1465 1265 1485 1285
rect 1465 1215 1485 1235
rect 1465 1165 1485 1185
rect 1465 1115 1485 1135
rect 1465 1065 1485 1085
rect 1465 1015 1485 1035
rect 1465 965 1485 985
rect 1465 915 1485 935
rect 1465 865 1485 885
rect 1465 815 1485 835
rect 1465 765 1485 785
rect 1465 715 1485 735
rect 1465 665 1485 685
rect 1465 615 1485 635
rect 1465 565 1485 585
rect 1465 515 1485 535
rect 1465 465 1485 485
rect 1465 415 1485 435
rect 1465 365 1485 385
rect 1465 315 1485 335
rect 1465 265 1485 285
rect 1465 215 1485 235
rect 1465 165 1485 185
rect 1765 2765 1785 2785
rect 1815 2765 1835 2785
rect 1865 2765 1885 2785
rect 1915 2765 1935 2785
rect 1965 2765 1985 2785
rect 2015 2765 2035 2785
rect 2065 2765 2085 2785
rect 2115 2765 2135 2785
rect 2165 2765 2185 2785
rect 2215 2765 2235 2785
rect 2265 2765 2285 2785
rect 2315 2765 2335 2785
rect 2365 2765 2385 2785
rect 2415 2765 2435 2785
rect 2465 2765 2485 2785
rect 2515 2765 2535 2785
rect 2565 2765 2585 2785
rect 2615 2765 2635 2785
rect 2665 2765 2685 2785
rect 2715 2765 2735 2785
rect 2765 2765 2785 2785
rect 1765 2715 1785 2735
rect 2765 2715 2785 2735
rect 1765 2665 1785 2685
rect 1765 2615 1785 2635
rect 1765 2565 1785 2585
rect 1765 2515 1785 2535
rect 1765 2465 1785 2485
rect 1765 2415 1785 2435
rect 1765 2365 1785 2385
rect 1765 2315 1785 2335
rect 1765 2265 1785 2285
rect 1765 2215 1785 2235
rect 1765 2165 1785 2185
rect 1765 2115 1785 2135
rect 1765 2065 1785 2085
rect 1765 2015 1785 2035
rect 2765 2665 2785 2685
rect 2765 2615 2785 2635
rect 2765 2565 2785 2585
rect 2765 2515 2785 2535
rect 2765 2465 2785 2485
rect 2765 2415 2785 2435
rect 2765 2365 2785 2385
rect 2765 2315 2785 2335
rect 2765 2265 2785 2285
rect 2765 2215 2785 2235
rect 2765 2165 2785 2185
rect 2765 2115 2785 2135
rect 2765 2065 2785 2085
rect 2765 2015 2785 2035
rect 1765 1965 1785 1985
rect 1765 1915 1785 1935
rect 1765 1865 1785 1885
rect 2765 1965 2785 1985
rect 2765 1915 2785 1935
rect 2765 1865 2785 1885
rect 1765 1815 1785 1835
rect 1765 1765 1785 1785
rect 1765 1715 1785 1735
rect 1765 1665 1785 1685
rect 1765 1615 1785 1635
rect 1765 1565 1785 1585
rect 1765 1515 1785 1535
rect 1765 1465 1785 1485
rect 1765 1415 1785 1435
rect 1765 1365 1785 1385
rect 1765 1315 1785 1335
rect 1765 1265 1785 1285
rect 1765 1215 1785 1235
rect 1765 1165 1785 1185
rect 2765 1815 2785 1835
rect 2765 1765 2785 1785
rect 2765 1715 2785 1735
rect 2765 1665 2785 1685
rect 2765 1615 2785 1635
rect 2765 1565 2785 1585
rect 2765 1515 2785 1535
rect 2765 1465 2785 1485
rect 2765 1415 2785 1435
rect 2765 1365 2785 1385
rect 2765 1315 2785 1335
rect 2765 1265 2785 1285
rect 2765 1215 2785 1235
rect 2765 1165 2785 1185
rect 1765 1115 1785 1135
rect 2765 1115 2785 1135
rect 1765 1065 1785 1085
rect 1815 1065 1835 1085
rect 1865 1065 1885 1085
rect 1915 1065 1935 1085
rect 1965 1065 1985 1085
rect 2015 1065 2035 1085
rect 2065 1065 2085 1085
rect 2115 1065 2135 1085
rect 2165 1065 2185 1085
rect 2215 1065 2235 1085
rect 2265 1065 2285 1085
rect 2315 1065 2335 1085
rect 2365 1065 2385 1085
rect 2415 1065 2435 1085
rect 2465 1065 2485 1085
rect 2515 1065 2535 1085
rect 2565 1065 2585 1085
rect 2615 1065 2635 1085
rect 2665 1065 2685 1085
rect 2715 1065 2735 1085
rect 2765 1065 2785 1085
rect 3065 3665 3085 3685
rect 3065 3615 3085 3635
rect 3065 3565 3085 3585
rect 3065 3515 3085 3535
rect 3065 3465 3085 3485
rect 3065 3415 3085 3435
rect 3065 3365 3085 3385
rect 3065 3315 3085 3335
rect 3065 3265 3085 3285
rect 3065 3215 3085 3235
rect 3065 3165 3085 3185
rect 3065 3115 3085 3135
rect 3065 3065 3085 3085
rect 3065 3015 3085 3035
rect 3065 2965 3085 2985
rect 3065 2915 3085 2935
rect 3065 2865 3085 2885
rect 3065 2815 3085 2835
rect 3065 2765 3085 2785
rect 3065 2715 3085 2735
rect 3065 2665 3085 2685
rect 3065 2615 3085 2635
rect 3065 2565 3085 2585
rect 3065 2515 3085 2535
rect 3065 2465 3085 2485
rect 3065 2415 3085 2435
rect 3065 2365 3085 2385
rect 3065 2315 3085 2335
rect 3065 2265 3085 2285
rect 3065 2215 3085 2235
rect 3065 2165 3085 2185
rect 3065 2115 3085 2135
rect 3065 2065 3085 2085
rect 3065 2015 3085 2035
rect 3065 1965 3085 1985
rect 3065 1915 3085 1935
rect 3065 1865 3085 1885
rect 3065 1815 3085 1835
rect 3065 1765 3085 1785
rect 3065 1715 3085 1735
rect 3065 1665 3085 1685
rect 3065 1615 3085 1635
rect 3065 1565 3085 1585
rect 3065 1515 3085 1535
rect 3065 1465 3085 1485
rect 3065 1415 3085 1435
rect 3065 1365 3085 1385
rect 3065 1315 3085 1335
rect 3065 1265 3085 1285
rect 3065 1215 3085 1235
rect 3065 1165 3085 1185
rect 3065 1115 3085 1135
rect 3065 1065 3085 1085
rect 3065 1015 3085 1035
rect 3065 965 3085 985
rect 3065 915 3085 935
rect 3065 865 3085 885
rect 3065 815 3085 835
rect 3065 765 3085 785
rect 3065 715 3085 735
rect 3065 665 3085 685
rect 3065 615 3085 635
rect 3065 565 3085 585
rect 3065 515 3085 535
rect 3065 465 3085 485
rect 3065 415 3085 435
rect 3065 365 3085 385
rect 3065 315 3085 335
rect 3065 265 3085 285
rect 3065 215 3085 235
rect 3065 165 3085 185
rect 1465 115 1485 135
rect 1465 65 1485 85
rect 3065 115 3085 135
rect 3065 65 3085 85
rect 1465 15 1485 35
rect 1515 15 1535 35
rect 1565 15 1585 35
rect 1615 15 1635 35
rect 1665 15 1685 35
rect 1715 15 1735 35
rect 1765 15 1785 35
rect 1815 15 1835 35
rect 1865 15 1885 35
rect 1915 15 1935 35
rect 1965 15 1985 35
rect 2015 15 2035 35
rect 2065 15 2085 35
rect 2115 15 2135 35
rect 2165 15 2185 35
rect 2215 15 2235 35
rect 2265 15 2285 35
rect 2315 15 2335 35
rect 2365 15 2385 35
rect 2415 15 2435 35
rect 2465 15 2485 35
rect 2515 15 2535 35
rect 2565 15 2585 35
rect 2615 15 2635 35
rect 2665 15 2685 35
rect 2715 15 2735 35
rect 2765 15 2785 35
rect 2815 15 2835 35
rect 2865 15 2885 35
rect 2915 15 2935 35
rect 2965 15 2985 35
rect 3015 15 3035 35
rect 3065 15 3085 35
<< nsubdiffcont >>
rect 1615 3665 1635 3685
rect 1665 3665 1685 3685
rect 1715 3665 1735 3685
rect 1765 3665 1785 3685
rect 1815 3665 1835 3685
rect 1865 3665 1885 3685
rect 1915 3665 1935 3685
rect 1965 3665 1985 3685
rect 2015 3665 2035 3685
rect 2065 3665 2085 3685
rect 2115 3665 2135 3685
rect 2165 3665 2185 3685
rect 2215 3665 2235 3685
rect 2265 3665 2285 3685
rect 2315 3665 2335 3685
rect 2365 3665 2385 3685
rect 2415 3665 2435 3685
rect 2465 3665 2485 3685
rect 2515 3665 2535 3685
rect 2565 3665 2585 3685
rect 2615 3665 2635 3685
rect 2665 3665 2685 3685
rect 2715 3665 2735 3685
rect 2765 3665 2785 3685
rect 2815 3665 2835 3685
rect 2865 3665 2885 3685
rect 2915 3665 2935 3685
rect 1615 3615 1635 3635
rect 2915 3615 2935 3635
rect 1615 3565 1635 3585
rect 1615 3515 1635 3535
rect 1615 3465 1635 3485
rect 1615 3415 1635 3435
rect 1615 3365 1635 3385
rect 1615 3315 1635 3335
rect 1615 3265 1635 3285
rect 1615 3215 1635 3235
rect 1615 3165 1635 3185
rect 1615 3115 1635 3135
rect 2915 3565 2935 3585
rect 2915 3515 2935 3535
rect 2915 3465 2935 3485
rect 2915 3415 2935 3435
rect 2915 3365 2935 3385
rect 2915 3315 2935 3335
rect 2915 3265 2935 3285
rect 2915 3215 2935 3235
rect 2915 3165 2935 3185
rect 2915 3115 2935 3135
rect 1615 3065 1635 3085
rect 1615 3015 1635 3035
rect 2915 3065 2935 3085
rect 2915 3015 2935 3035
rect 1615 2965 1635 2985
rect 2915 2965 2935 2985
rect 1615 2915 1635 2935
rect 1665 2915 1685 2935
rect 1715 2915 1735 2935
rect 1765 2915 1785 2935
rect 1815 2915 1835 2935
rect 1865 2915 1885 2935
rect 1915 2915 1935 2935
rect 1965 2915 1985 2935
rect 2015 2915 2035 2935
rect 2065 2915 2085 2935
rect 2115 2915 2135 2935
rect 2165 2915 2185 2935
rect 2215 2915 2235 2935
rect 2265 2915 2285 2935
rect 2315 2915 2335 2935
rect 2365 2915 2385 2935
rect 2415 2915 2435 2935
rect 2465 2915 2485 2935
rect 2515 2915 2535 2935
rect 2565 2915 2585 2935
rect 2615 2915 2635 2935
rect 2665 2915 2685 2935
rect 2715 2915 2735 2935
rect 2765 2915 2785 2935
rect 2815 2915 2835 2935
rect 2865 2915 2885 2935
rect 2915 2915 2935 2935
rect 1615 2865 1635 2885
rect 1615 2815 1635 2835
rect 2915 2865 2935 2885
rect 2915 2815 2935 2835
rect 1615 2765 1635 2785
rect 1615 2715 1635 2735
rect 1615 2665 1635 2685
rect 1615 2615 1635 2635
rect 1615 2565 1635 2585
rect 1615 2515 1635 2535
rect 1615 2465 1635 2485
rect 1615 2415 1635 2435
rect 1615 2365 1635 2385
rect 1615 2315 1635 2335
rect 1615 2265 1635 2285
rect 1615 2215 1635 2235
rect 1615 2165 1635 2185
rect 1615 2115 1635 2135
rect 1615 2065 1635 2085
rect 1615 2015 1635 2035
rect 1615 1965 1635 1985
rect 1615 1915 1635 1935
rect 1615 1865 1635 1885
rect 1615 1815 1635 1835
rect 1615 1765 1635 1785
rect 1615 1715 1635 1735
rect 1615 1665 1635 1685
rect 1615 1615 1635 1635
rect 1615 1565 1635 1585
rect 1615 1515 1635 1535
rect 1615 1465 1635 1485
rect 1615 1415 1635 1435
rect 1615 1365 1635 1385
rect 1615 1315 1635 1335
rect 1615 1265 1635 1285
rect 1615 1215 1635 1235
rect 1615 1165 1635 1185
rect 1615 1115 1635 1135
rect 1615 1065 1635 1085
rect 2915 2765 2935 2785
rect 2915 2715 2935 2735
rect 2915 2665 2935 2685
rect 2915 2615 2935 2635
rect 2915 2565 2935 2585
rect 2915 2515 2935 2535
rect 2915 2465 2935 2485
rect 2915 2415 2935 2435
rect 2915 2365 2935 2385
rect 2915 2315 2935 2335
rect 2915 2265 2935 2285
rect 2915 2215 2935 2235
rect 2915 2165 2935 2185
rect 2915 2115 2935 2135
rect 2915 2065 2935 2085
rect 2915 2015 2935 2035
rect 2915 1965 2935 1985
rect 2915 1915 2935 1935
rect 2915 1865 2935 1885
rect 2915 1815 2935 1835
rect 2915 1765 2935 1785
rect 2915 1715 2935 1735
rect 2915 1665 2935 1685
rect 2915 1615 2935 1635
rect 2915 1565 2935 1585
rect 2915 1515 2935 1535
rect 2915 1465 2935 1485
rect 2915 1415 2935 1435
rect 2915 1365 2935 1385
rect 2915 1315 2935 1335
rect 2915 1265 2935 1285
rect 2915 1215 2935 1235
rect 2915 1165 2935 1185
rect 2915 1115 2935 1135
rect 2915 1065 2935 1085
rect 1615 1015 1635 1035
rect 1615 965 1635 985
rect 2915 1015 2935 1035
rect 2915 965 2935 985
rect 1615 915 1635 935
rect 1665 915 1685 935
rect 1715 915 1735 935
rect 1765 915 1785 935
rect 1815 915 1835 935
rect 1865 915 1885 935
rect 1915 915 1935 935
rect 1965 915 1985 935
rect 2015 915 2035 935
rect 2065 915 2085 935
rect 2115 915 2135 935
rect 2165 915 2185 935
rect 2215 915 2235 935
rect 2265 915 2285 935
rect 2315 915 2335 935
rect 2365 915 2385 935
rect 2415 915 2435 935
rect 2465 915 2485 935
rect 2515 915 2535 935
rect 2565 915 2585 935
rect 2615 915 2635 935
rect 2665 915 2685 935
rect 2715 915 2735 935
rect 2765 915 2785 935
rect 2815 915 2835 935
rect 2865 915 2885 935
rect 2915 915 2935 935
rect 1615 865 1635 885
rect 2915 865 2935 885
rect 1615 815 1635 835
rect 1615 765 1635 785
rect 2915 815 2935 835
rect 2915 765 2935 785
rect 1615 715 1635 735
rect 1615 665 1635 685
rect 1615 615 1635 635
rect 1615 565 1635 585
rect 1615 515 1635 535
rect 1615 465 1635 485
rect 1615 415 1635 435
rect 1615 365 1635 385
rect 1615 315 1635 335
rect 1615 265 1635 285
rect 2915 715 2935 735
rect 2915 665 2935 685
rect 2915 615 2935 635
rect 2915 565 2935 585
rect 2915 515 2935 535
rect 2915 465 2935 485
rect 2915 415 2935 435
rect 2915 365 2935 385
rect 2915 315 2935 335
rect 2915 265 2935 285
rect 1615 215 1635 235
rect 2915 215 2935 235
rect 1615 165 1635 185
rect 1665 165 1685 185
rect 1715 165 1735 185
rect 1765 165 1785 185
rect 1815 165 1835 185
rect 1865 165 1885 185
rect 1915 165 1935 185
rect 1965 165 1985 185
rect 2015 165 2035 185
rect 2065 165 2085 185
rect 2115 165 2135 185
rect 2165 165 2185 185
rect 2215 165 2235 185
rect 2265 165 2285 185
rect 2315 165 2335 185
rect 2365 165 2385 185
rect 2415 165 2435 185
rect 2465 165 2485 185
rect 2515 165 2535 185
rect 2565 165 2585 185
rect 2615 165 2635 185
rect 2665 165 2685 185
rect 2715 165 2735 185
rect 2765 165 2785 185
rect 2815 165 2835 185
rect 2865 165 2885 185
rect 2915 165 2935 185
<< poly >>
rect 1900 3600 1950 3615
rect 2000 3600 2050 3615
rect 2100 3600 2150 3615
rect 2200 3600 2250 3615
rect 2300 3600 2350 3615
rect 2400 3600 2450 3615
rect 2500 3600 2550 3615
rect 2600 3600 2650 3615
rect 1900 3050 1950 3100
rect 2000 3050 2050 3100
rect 1900 3035 2050 3050
rect 1900 3015 1915 3035
rect 1935 3015 1965 3035
rect 1985 3015 2015 3035
rect 2035 3015 2050 3035
rect 1900 3000 2050 3015
rect 2100 3050 2150 3100
rect 2200 3050 2250 3100
rect 2100 3035 2250 3050
rect 2100 3015 2115 3035
rect 2135 3015 2165 3035
rect 2185 3015 2215 3035
rect 2235 3015 2250 3035
rect 2100 3000 2250 3015
rect 2300 3050 2350 3100
rect 2400 3050 2450 3100
rect 2300 3035 2450 3050
rect 2300 3015 2315 3035
rect 2335 3015 2365 3035
rect 2385 3015 2415 3035
rect 2435 3015 2450 3035
rect 2300 3000 2450 3015
rect 2500 3050 2550 3100
rect 2600 3050 2650 3100
rect 2500 3035 2650 3050
rect 2500 3015 2515 3035
rect 2535 3015 2565 3035
rect 2585 3015 2615 3035
rect 2635 3015 2650 3035
rect 2500 3000 2650 3015
rect 1900 2700 1950 2715
rect 2000 2700 2050 2715
rect 2100 2700 2150 2715
rect 2200 2700 2250 2715
rect 2300 2700 2350 2715
rect 2400 2700 2450 2715
rect 2500 2700 2550 2715
rect 2600 2700 2650 2715
rect 1900 1950 1950 2000
rect 2000 1950 2050 2000
rect 1900 1935 2050 1950
rect 1900 1915 1915 1935
rect 1935 1915 1965 1935
rect 1985 1915 2015 1935
rect 2035 1915 2050 1935
rect 1900 1900 2050 1915
rect 1900 1850 1950 1900
rect 2000 1850 2050 1900
rect 2100 1950 2150 2000
rect 2200 1950 2250 2000
rect 2100 1935 2250 1950
rect 2100 1915 2115 1935
rect 2135 1915 2165 1935
rect 2185 1915 2215 1935
rect 2235 1915 2250 1935
rect 2100 1900 2250 1915
rect 2100 1850 2150 1900
rect 2200 1850 2250 1900
rect 2300 1950 2350 2000
rect 2400 1950 2450 2000
rect 2300 1935 2450 1950
rect 2300 1915 2315 1935
rect 2335 1915 2365 1935
rect 2385 1915 2415 1935
rect 2435 1915 2450 1935
rect 2300 1900 2450 1915
rect 2300 1850 2350 1900
rect 2400 1850 2450 1900
rect 2500 1950 2550 2000
rect 2600 1950 2650 2000
rect 2500 1935 2650 1950
rect 2500 1915 2515 1935
rect 2535 1915 2565 1935
rect 2585 1915 2615 1935
rect 2635 1915 2650 1935
rect 2500 1900 2650 1915
rect 2500 1850 2550 1900
rect 2600 1850 2650 1900
rect 1900 1135 1950 1150
rect 2000 1135 2050 1150
rect 2100 1135 2150 1150
rect 2200 1135 2250 1150
rect 2300 1135 2350 1150
rect 2400 1135 2450 1150
rect 2500 1135 2550 1150
rect 2600 1135 2650 1150
rect 1900 835 2050 850
rect 1900 815 1915 835
rect 1935 815 1965 835
rect 1985 815 2015 835
rect 2035 815 2050 835
rect 1900 800 2050 815
rect 1900 750 1950 800
rect 2000 750 2050 800
rect 2100 835 2250 850
rect 2100 815 2115 835
rect 2135 815 2165 835
rect 2185 815 2215 835
rect 2235 815 2250 835
rect 2100 800 2250 815
rect 2100 750 2150 800
rect 2200 750 2250 800
rect 2300 835 2450 850
rect 2300 815 2315 835
rect 2335 815 2365 835
rect 2385 815 2415 835
rect 2435 815 2450 835
rect 2300 800 2450 815
rect 2300 750 2350 800
rect 2400 750 2450 800
rect 2500 835 2650 850
rect 2500 815 2515 835
rect 2535 815 2565 835
rect 2585 815 2615 835
rect 2635 815 2650 835
rect 2500 800 2650 815
rect 2500 750 2550 800
rect 2600 750 2650 800
rect 1900 235 1950 250
rect 2000 235 2050 250
rect 2100 235 2150 250
rect 2200 235 2250 250
rect 2300 235 2350 250
rect 2400 235 2450 250
rect 2500 235 2550 250
rect 2600 235 2650 250
<< polycont >>
rect 1915 3015 1935 3035
rect 1965 3015 1985 3035
rect 2015 3015 2035 3035
rect 2115 3015 2135 3035
rect 2165 3015 2185 3035
rect 2215 3015 2235 3035
rect 2315 3015 2335 3035
rect 2365 3015 2385 3035
rect 2415 3015 2435 3035
rect 2515 3015 2535 3035
rect 2565 3015 2585 3035
rect 2615 3015 2635 3035
rect 1915 1915 1935 1935
rect 1965 1915 1985 1935
rect 2015 1915 2035 1935
rect 2115 1915 2135 1935
rect 2165 1915 2185 1935
rect 2215 1915 2235 1935
rect 2315 1915 2335 1935
rect 2365 1915 2385 1935
rect 2415 1915 2435 1935
rect 2515 1915 2535 1935
rect 2565 1915 2585 1935
rect 2615 1915 2635 1935
rect 1915 815 1935 835
rect 1965 815 1985 835
rect 2015 815 2035 835
rect 2115 815 2135 835
rect 2165 815 2185 835
rect 2215 815 2235 835
rect 2315 815 2335 835
rect 2365 815 2385 835
rect 2415 815 2435 835
rect 2515 815 2535 835
rect 2565 815 2585 835
rect 2615 815 2635 835
<< locali >>
rect 1450 3835 3100 3850
rect 1450 3815 1465 3835
rect 1485 3815 1515 3835
rect 1535 3815 1565 3835
rect 1585 3815 1615 3835
rect 1635 3815 1665 3835
rect 1685 3815 1715 3835
rect 1735 3815 1765 3835
rect 1785 3815 1815 3835
rect 1835 3815 1865 3835
rect 1885 3815 1915 3835
rect 1935 3815 1965 3835
rect 1985 3815 2015 3835
rect 2035 3815 2065 3835
rect 2085 3815 2115 3835
rect 2135 3815 2165 3835
rect 2185 3815 2215 3835
rect 2235 3815 2265 3835
rect 2285 3815 2315 3835
rect 2335 3815 2365 3835
rect 2385 3815 2415 3835
rect 2435 3815 2465 3835
rect 2485 3815 2515 3835
rect 2535 3815 2565 3835
rect 2585 3815 2615 3835
rect 2635 3815 2665 3835
rect 2685 3815 2715 3835
rect 2735 3815 2765 3835
rect 2785 3815 2815 3835
rect 2835 3815 2865 3835
rect 2885 3815 2915 3835
rect 2935 3815 2965 3835
rect 2985 3815 3015 3835
rect 3035 3815 3065 3835
rect 3085 3815 3100 3835
rect 1450 3800 3100 3815
rect 1450 3785 1500 3800
rect 1450 3765 1465 3785
rect 1485 3765 1500 3785
rect 1450 3735 1500 3765
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1450 3685 1500 3715
rect 3050 3785 3100 3800
rect 3050 3765 3065 3785
rect 3085 3765 3100 3785
rect 3050 3735 3100 3765
rect 3050 3715 3065 3735
rect 3085 3715 3100 3735
rect 1450 3665 1465 3685
rect 1485 3665 1500 3685
rect 1450 3635 1500 3665
rect 1450 3615 1465 3635
rect 1485 3615 1500 3635
rect 1450 3585 1500 3615
rect 1450 3565 1465 3585
rect 1485 3565 1500 3585
rect 1450 3535 1500 3565
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3285 1500 3315
rect 1450 3265 1465 3285
rect 1485 3265 1500 3285
rect 1450 3235 1500 3265
rect 1450 3215 1465 3235
rect 1485 3215 1500 3235
rect 1450 3185 1500 3215
rect 1450 3165 1465 3185
rect 1485 3165 1500 3185
rect 1450 3135 1500 3165
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3085 1500 3115
rect 1450 3065 1465 3085
rect 1485 3065 1500 3085
rect 1450 3035 1500 3065
rect 1450 3015 1465 3035
rect 1485 3015 1500 3035
rect 1450 2985 1500 3015
rect 1450 2965 1465 2985
rect 1485 2965 1500 2985
rect 1450 2935 1500 2965
rect 1450 2915 1465 2935
rect 1485 2915 1500 2935
rect 1450 2885 1500 2915
rect 1450 2865 1465 2885
rect 1485 2865 1500 2885
rect 1450 2835 1500 2865
rect 1450 2815 1465 2835
rect 1485 2815 1500 2835
rect 1450 2785 1500 2815
rect 1450 2765 1465 2785
rect 1485 2765 1500 2785
rect 1450 2735 1500 2765
rect 1450 2715 1465 2735
rect 1485 2715 1500 2735
rect 1450 2685 1500 2715
rect 1450 2665 1465 2685
rect 1485 2665 1500 2685
rect 1450 2635 1500 2665
rect 1450 2615 1465 2635
rect 1485 2615 1500 2635
rect 1450 2585 1500 2615
rect 1450 2565 1465 2585
rect 1485 2565 1500 2585
rect 1450 2535 1500 2565
rect 1450 2515 1465 2535
rect 1485 2515 1500 2535
rect 1450 2485 1500 2515
rect 1450 2465 1465 2485
rect 1485 2465 1500 2485
rect 1450 2435 1500 2465
rect 1450 2415 1465 2435
rect 1485 2415 1500 2435
rect 1450 2385 1500 2415
rect 1450 2365 1465 2385
rect 1485 2365 1500 2385
rect 1450 2335 1500 2365
rect 1450 2315 1465 2335
rect 1485 2315 1500 2335
rect 1450 2285 1500 2315
rect 1450 2265 1465 2285
rect 1485 2265 1500 2285
rect 1450 2235 1500 2265
rect 1450 2215 1465 2235
rect 1485 2215 1500 2235
rect 1450 2185 1500 2215
rect 1450 2165 1465 2185
rect 1485 2165 1500 2185
rect 1450 2135 1500 2165
rect 1450 2115 1465 2135
rect 1485 2115 1500 2135
rect 1450 2085 1500 2115
rect 1450 2065 1465 2085
rect 1485 2065 1500 2085
rect 1450 2035 1500 2065
rect 1450 2015 1465 2035
rect 1485 2015 1500 2035
rect 1450 1985 1500 2015
rect 1450 1965 1465 1985
rect 1485 1965 1500 1985
rect 1450 1935 1500 1965
rect 1450 1915 1465 1935
rect 1485 1915 1500 1935
rect 1450 1885 1500 1915
rect 1450 1865 1465 1885
rect 1485 1865 1500 1885
rect 1450 1835 1500 1865
rect 1450 1815 1465 1835
rect 1485 1815 1500 1835
rect 1450 1785 1500 1815
rect 1450 1765 1465 1785
rect 1485 1765 1500 1785
rect 1450 1735 1500 1765
rect 1450 1715 1465 1735
rect 1485 1715 1500 1735
rect 1450 1685 1500 1715
rect 1450 1665 1465 1685
rect 1485 1665 1500 1685
rect 1450 1635 1500 1665
rect 1450 1615 1465 1635
rect 1485 1615 1500 1635
rect 1450 1585 1500 1615
rect 1450 1565 1465 1585
rect 1485 1565 1500 1585
rect 1450 1535 1500 1565
rect 1450 1515 1465 1535
rect 1485 1515 1500 1535
rect 1450 1485 1500 1515
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 935 1500 965
rect 1450 915 1465 935
rect 1485 915 1500 935
rect 1450 885 1500 915
rect 1450 865 1465 885
rect 1485 865 1500 885
rect 1450 835 1500 865
rect 1450 815 1465 835
rect 1485 815 1500 835
rect 1450 785 1500 815
rect 1450 765 1465 785
rect 1485 765 1500 785
rect 1450 735 1500 765
rect 1450 715 1465 735
rect 1485 715 1500 735
rect 1450 685 1500 715
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 135 1500 165
rect 1600 3685 2950 3700
rect 1600 3665 1615 3685
rect 1635 3665 1665 3685
rect 1685 3665 1715 3685
rect 1735 3665 1765 3685
rect 1785 3665 1815 3685
rect 1835 3665 1865 3685
rect 1885 3665 1915 3685
rect 1935 3665 1965 3685
rect 1985 3665 2015 3685
rect 2035 3665 2065 3685
rect 2085 3665 2115 3685
rect 2135 3665 2165 3685
rect 2185 3665 2215 3685
rect 2235 3665 2265 3685
rect 2285 3665 2315 3685
rect 2335 3665 2365 3685
rect 2385 3665 2415 3685
rect 2435 3665 2465 3685
rect 2485 3665 2515 3685
rect 2535 3665 2565 3685
rect 2585 3665 2615 3685
rect 2635 3665 2665 3685
rect 2685 3665 2715 3685
rect 2735 3665 2765 3685
rect 2785 3665 2815 3685
rect 2835 3665 2865 3685
rect 2885 3665 2915 3685
rect 2935 3665 2950 3685
rect 1600 3650 2950 3665
rect 1600 3635 1650 3650
rect 1600 3615 1615 3635
rect 1635 3615 1650 3635
rect 1600 3585 1650 3615
rect 1600 3565 1615 3585
rect 1635 3565 1650 3585
rect 1600 3535 1650 3565
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3285 1650 3315
rect 1600 3265 1615 3285
rect 1635 3265 1650 3285
rect 1600 3235 1650 3265
rect 1600 3215 1615 3235
rect 1635 3215 1650 3235
rect 1600 3185 1650 3215
rect 1600 3165 1615 3185
rect 1635 3165 1650 3185
rect 1600 3135 1650 3165
rect 1600 3115 1615 3135
rect 1635 3115 1650 3135
rect 1600 3085 1650 3115
rect 1850 3585 1900 3600
rect 1850 3565 1865 3585
rect 1885 3565 1900 3585
rect 1850 3535 1900 3565
rect 1850 3515 1865 3535
rect 1885 3515 1900 3535
rect 1850 3485 1900 3515
rect 1850 3465 1865 3485
rect 1885 3465 1900 3485
rect 1850 3435 1900 3465
rect 1850 3415 1865 3435
rect 1885 3415 1900 3435
rect 1850 3385 1900 3415
rect 1850 3365 1865 3385
rect 1885 3365 1900 3385
rect 1850 3335 1900 3365
rect 1850 3315 1865 3335
rect 1885 3315 1900 3335
rect 1850 3285 1900 3315
rect 1850 3265 1865 3285
rect 1885 3265 1900 3285
rect 1850 3235 1900 3265
rect 1850 3215 1865 3235
rect 1885 3215 1900 3235
rect 1850 3185 1900 3215
rect 1850 3165 1865 3185
rect 1885 3165 1900 3185
rect 1850 3135 1900 3165
rect 1850 3115 1865 3135
rect 1885 3115 1900 3135
rect 1850 3100 1900 3115
rect 1950 3585 2000 3600
rect 1950 3565 1965 3585
rect 1985 3565 2000 3585
rect 1950 3535 2000 3565
rect 1950 3515 1965 3535
rect 1985 3515 2000 3535
rect 1950 3485 2000 3515
rect 1950 3465 1965 3485
rect 1985 3465 2000 3485
rect 1950 3435 2000 3465
rect 1950 3415 1965 3435
rect 1985 3415 2000 3435
rect 1950 3385 2000 3415
rect 1950 3365 1965 3385
rect 1985 3365 2000 3385
rect 1950 3335 2000 3365
rect 1950 3315 1965 3335
rect 1985 3315 2000 3335
rect 1950 3285 2000 3315
rect 1950 3265 1965 3285
rect 1985 3265 2000 3285
rect 1950 3235 2000 3265
rect 1950 3215 1965 3235
rect 1985 3215 2000 3235
rect 1950 3185 2000 3215
rect 1950 3165 1965 3185
rect 1985 3165 2000 3185
rect 1950 3135 2000 3165
rect 1950 3115 1965 3135
rect 1985 3115 2000 3135
rect 1950 3100 2000 3115
rect 2050 3585 2100 3600
rect 2050 3565 2065 3585
rect 2085 3565 2100 3585
rect 2050 3535 2100 3565
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3285 2100 3315
rect 2050 3265 2065 3285
rect 2085 3265 2100 3285
rect 2050 3235 2100 3265
rect 2050 3215 2065 3235
rect 2085 3215 2100 3235
rect 2050 3185 2100 3215
rect 2050 3165 2065 3185
rect 2085 3165 2100 3185
rect 2050 3135 2100 3165
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3100 2100 3115
rect 2150 3585 2200 3600
rect 2150 3565 2165 3585
rect 2185 3565 2200 3585
rect 2150 3535 2200 3565
rect 2150 3515 2165 3535
rect 2185 3515 2200 3535
rect 2150 3485 2200 3515
rect 2150 3465 2165 3485
rect 2185 3465 2200 3485
rect 2150 3435 2200 3465
rect 2150 3415 2165 3435
rect 2185 3415 2200 3435
rect 2150 3385 2200 3415
rect 2150 3365 2165 3385
rect 2185 3365 2200 3385
rect 2150 3335 2200 3365
rect 2150 3315 2165 3335
rect 2185 3315 2200 3335
rect 2150 3285 2200 3315
rect 2150 3265 2165 3285
rect 2185 3265 2200 3285
rect 2150 3235 2200 3265
rect 2150 3215 2165 3235
rect 2185 3215 2200 3235
rect 2150 3185 2200 3215
rect 2150 3165 2165 3185
rect 2185 3165 2200 3185
rect 2150 3135 2200 3165
rect 2150 3115 2165 3135
rect 2185 3115 2200 3135
rect 2150 3100 2200 3115
rect 2250 3585 2300 3650
rect 2900 3635 2950 3650
rect 2900 3615 2915 3635
rect 2935 3615 2950 3635
rect 2250 3565 2265 3585
rect 2285 3565 2300 3585
rect 2250 3535 2300 3565
rect 2250 3515 2265 3535
rect 2285 3515 2300 3535
rect 2250 3485 2300 3515
rect 2250 3465 2265 3485
rect 2285 3465 2300 3485
rect 2250 3435 2300 3465
rect 2250 3415 2265 3435
rect 2285 3415 2300 3435
rect 2250 3385 2300 3415
rect 2250 3365 2265 3385
rect 2285 3365 2300 3385
rect 2250 3335 2300 3365
rect 2250 3315 2265 3335
rect 2285 3315 2300 3335
rect 2250 3285 2300 3315
rect 2250 3265 2265 3285
rect 2285 3265 2300 3285
rect 2250 3235 2300 3265
rect 2250 3215 2265 3235
rect 2285 3215 2300 3235
rect 2250 3185 2300 3215
rect 2250 3165 2265 3185
rect 2285 3165 2300 3185
rect 2250 3135 2300 3165
rect 2250 3115 2265 3135
rect 2285 3115 2300 3135
rect 2250 3100 2300 3115
rect 2350 3585 2400 3600
rect 2350 3565 2365 3585
rect 2385 3565 2400 3585
rect 2350 3535 2400 3565
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3285 2400 3315
rect 2350 3265 2365 3285
rect 2385 3265 2400 3285
rect 2350 3235 2400 3265
rect 2350 3215 2365 3235
rect 2385 3215 2400 3235
rect 2350 3185 2400 3215
rect 2350 3165 2365 3185
rect 2385 3165 2400 3185
rect 2350 3135 2400 3165
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3100 2400 3115
rect 2450 3585 2500 3600
rect 2450 3565 2465 3585
rect 2485 3565 2500 3585
rect 2450 3535 2500 3565
rect 2450 3515 2465 3535
rect 2485 3515 2500 3535
rect 2450 3485 2500 3515
rect 2450 3465 2465 3485
rect 2485 3465 2500 3485
rect 2450 3435 2500 3465
rect 2450 3415 2465 3435
rect 2485 3415 2500 3435
rect 2450 3385 2500 3415
rect 2450 3365 2465 3385
rect 2485 3365 2500 3385
rect 2450 3335 2500 3365
rect 2450 3315 2465 3335
rect 2485 3315 2500 3335
rect 2450 3285 2500 3315
rect 2450 3265 2465 3285
rect 2485 3265 2500 3285
rect 2450 3235 2500 3265
rect 2450 3215 2465 3235
rect 2485 3215 2500 3235
rect 2450 3185 2500 3215
rect 2450 3165 2465 3185
rect 2485 3165 2500 3185
rect 2450 3135 2500 3165
rect 2450 3115 2465 3135
rect 2485 3115 2500 3135
rect 2450 3100 2500 3115
rect 2550 3585 2600 3600
rect 2550 3565 2565 3585
rect 2585 3565 2600 3585
rect 2550 3535 2600 3565
rect 2550 3515 2565 3535
rect 2585 3515 2600 3535
rect 2550 3485 2600 3515
rect 2550 3465 2565 3485
rect 2585 3465 2600 3485
rect 2550 3435 2600 3465
rect 2550 3415 2565 3435
rect 2585 3415 2600 3435
rect 2550 3385 2600 3415
rect 2550 3365 2565 3385
rect 2585 3365 2600 3385
rect 2550 3335 2600 3365
rect 2550 3315 2565 3335
rect 2585 3315 2600 3335
rect 2550 3285 2600 3315
rect 2550 3265 2565 3285
rect 2585 3265 2600 3285
rect 2550 3235 2600 3265
rect 2550 3215 2565 3235
rect 2585 3215 2600 3235
rect 2550 3185 2600 3215
rect 2550 3165 2565 3185
rect 2585 3165 2600 3185
rect 2550 3135 2600 3165
rect 2550 3115 2565 3135
rect 2585 3115 2600 3135
rect 2550 3100 2600 3115
rect 2650 3585 2700 3600
rect 2650 3565 2665 3585
rect 2685 3565 2700 3585
rect 2650 3535 2700 3565
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3285 2700 3315
rect 2650 3265 2665 3285
rect 2685 3265 2700 3285
rect 2650 3235 2700 3265
rect 2650 3215 2665 3235
rect 2685 3215 2700 3235
rect 2650 3185 2700 3215
rect 2650 3165 2665 3185
rect 2685 3165 2700 3185
rect 2650 3135 2700 3165
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3100 2700 3115
rect 2900 3585 2950 3615
rect 2900 3565 2915 3585
rect 2935 3565 2950 3585
rect 2900 3535 2950 3565
rect 2900 3515 2915 3535
rect 2935 3515 2950 3535
rect 2900 3485 2950 3515
rect 2900 3465 2915 3485
rect 2935 3465 2950 3485
rect 2900 3435 2950 3465
rect 2900 3415 2915 3435
rect 2935 3415 2950 3435
rect 2900 3385 2950 3415
rect 2900 3365 2915 3385
rect 2935 3365 2950 3385
rect 2900 3335 2950 3365
rect 2900 3315 2915 3335
rect 2935 3315 2950 3335
rect 2900 3285 2950 3315
rect 2900 3265 2915 3285
rect 2935 3265 2950 3285
rect 2900 3235 2950 3265
rect 2900 3215 2915 3235
rect 2935 3215 2950 3235
rect 2900 3185 2950 3215
rect 2900 3165 2915 3185
rect 2935 3165 2950 3185
rect 2900 3135 2950 3165
rect 2900 3115 2915 3135
rect 2935 3115 2950 3135
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1600 3035 1650 3065
rect 2900 3085 2950 3115
rect 2900 3065 2915 3085
rect 2935 3065 2950 3085
rect 1600 3015 1615 3035
rect 1635 3015 1650 3035
rect 1600 2985 1650 3015
rect 1900 3035 2050 3050
rect 1900 3015 1915 3035
rect 1935 3015 1965 3035
rect 1985 3015 2015 3035
rect 2035 3015 2050 3035
rect 1900 3000 2050 3015
rect 2100 3035 2250 3050
rect 2100 3015 2115 3035
rect 2135 3015 2165 3035
rect 2185 3015 2215 3035
rect 2235 3015 2250 3035
rect 2100 3000 2250 3015
rect 2300 3035 2450 3050
rect 2300 3015 2315 3035
rect 2335 3015 2365 3035
rect 2385 3015 2415 3035
rect 2435 3015 2450 3035
rect 2300 3000 2450 3015
rect 2500 3035 2650 3050
rect 2500 3015 2515 3035
rect 2535 3015 2565 3035
rect 2585 3015 2615 3035
rect 2635 3015 2650 3035
rect 2500 3000 2650 3015
rect 2900 3035 2950 3065
rect 2900 3015 2915 3035
rect 2935 3015 2950 3035
rect 1600 2965 1615 2985
rect 1635 2965 1650 2985
rect 1600 2950 1650 2965
rect 2900 2985 2950 3015
rect 2900 2965 2915 2985
rect 2935 2965 2950 2985
rect 2900 2950 2950 2965
rect 1600 2935 2950 2950
rect 1600 2915 1615 2935
rect 1635 2915 1665 2935
rect 1685 2915 1715 2935
rect 1735 2915 1765 2935
rect 1785 2915 1815 2935
rect 1835 2915 1865 2935
rect 1885 2915 1915 2935
rect 1935 2915 1965 2935
rect 1985 2915 2015 2935
rect 2035 2915 2065 2935
rect 2085 2915 2115 2935
rect 2135 2915 2165 2935
rect 2185 2915 2215 2935
rect 2235 2915 2265 2935
rect 2285 2915 2315 2935
rect 2335 2915 2365 2935
rect 2385 2915 2415 2935
rect 2435 2915 2465 2935
rect 2485 2915 2515 2935
rect 2535 2915 2565 2935
rect 2585 2915 2615 2935
rect 2635 2915 2665 2935
rect 2685 2915 2715 2935
rect 2735 2915 2765 2935
rect 2785 2915 2815 2935
rect 2835 2915 2865 2935
rect 2885 2915 2915 2935
rect 2935 2915 2950 2935
rect 1600 2900 2950 2915
rect 1600 2885 1650 2900
rect 1600 2865 1615 2885
rect 1635 2865 1650 2885
rect 1600 2835 1650 2865
rect 1600 2815 1615 2835
rect 1635 2815 1650 2835
rect 1600 2785 1650 2815
rect 2900 2885 2950 2900
rect 2900 2865 2915 2885
rect 2935 2865 2950 2885
rect 2900 2835 2950 2865
rect 2900 2815 2915 2835
rect 2935 2815 2950 2835
rect 1600 2765 1615 2785
rect 1635 2765 1650 2785
rect 1600 2735 1650 2765
rect 1600 2715 1615 2735
rect 1635 2715 1650 2735
rect 1600 2685 1650 2715
rect 1600 2665 1615 2685
rect 1635 2665 1650 2685
rect 1600 2635 1650 2665
rect 1600 2615 1615 2635
rect 1635 2615 1650 2635
rect 1600 2585 1650 2615
rect 1600 2565 1615 2585
rect 1635 2565 1650 2585
rect 1600 2535 1650 2565
rect 1600 2515 1615 2535
rect 1635 2515 1650 2535
rect 1600 2485 1650 2515
rect 1600 2465 1615 2485
rect 1635 2465 1650 2485
rect 1600 2435 1650 2465
rect 1600 2415 1615 2435
rect 1635 2415 1650 2435
rect 1600 2385 1650 2415
rect 1600 2365 1615 2385
rect 1635 2365 1650 2385
rect 1600 2335 1650 2365
rect 1600 2315 1615 2335
rect 1635 2315 1650 2335
rect 1600 2285 1650 2315
rect 1600 2265 1615 2285
rect 1635 2265 1650 2285
rect 1600 2235 1650 2265
rect 1600 2215 1615 2235
rect 1635 2215 1650 2235
rect 1600 2185 1650 2215
rect 1600 2165 1615 2185
rect 1635 2165 1650 2185
rect 1600 2135 1650 2165
rect 1600 2115 1615 2135
rect 1635 2115 1650 2135
rect 1600 2085 1650 2115
rect 1600 2065 1615 2085
rect 1635 2065 1650 2085
rect 1600 2035 1650 2065
rect 1600 2015 1615 2035
rect 1635 2015 1650 2035
rect 1600 1985 1650 2015
rect 1600 1965 1615 1985
rect 1635 1965 1650 1985
rect 1600 1935 1650 1965
rect 1600 1915 1615 1935
rect 1635 1915 1650 1935
rect 1600 1885 1650 1915
rect 1600 1865 1615 1885
rect 1635 1865 1650 1885
rect 1600 1835 1650 1865
rect 1600 1815 1615 1835
rect 1635 1815 1650 1835
rect 1600 1785 1650 1815
rect 1600 1765 1615 1785
rect 1635 1765 1650 1785
rect 1600 1735 1650 1765
rect 1600 1715 1615 1735
rect 1635 1715 1650 1735
rect 1600 1685 1650 1715
rect 1600 1665 1615 1685
rect 1635 1665 1650 1685
rect 1600 1635 1650 1665
rect 1600 1615 1615 1635
rect 1635 1615 1650 1635
rect 1600 1585 1650 1615
rect 1600 1565 1615 1585
rect 1635 1565 1650 1585
rect 1600 1535 1650 1565
rect 1600 1515 1615 1535
rect 1635 1515 1650 1535
rect 1600 1485 1650 1515
rect 1600 1465 1615 1485
rect 1635 1465 1650 1485
rect 1600 1435 1650 1465
rect 1600 1415 1615 1435
rect 1635 1415 1650 1435
rect 1600 1385 1650 1415
rect 1600 1365 1615 1385
rect 1635 1365 1650 1385
rect 1600 1335 1650 1365
rect 1600 1315 1615 1335
rect 1635 1315 1650 1335
rect 1600 1285 1650 1315
rect 1600 1265 1615 1285
rect 1635 1265 1650 1285
rect 1600 1235 1650 1265
rect 1600 1215 1615 1235
rect 1635 1215 1650 1235
rect 1600 1185 1650 1215
rect 1600 1165 1615 1185
rect 1635 1165 1650 1185
rect 1600 1135 1650 1165
rect 1600 1115 1615 1135
rect 1635 1115 1650 1135
rect 1600 1085 1650 1115
rect 1600 1065 1615 1085
rect 1635 1065 1650 1085
rect 1600 1035 1650 1065
rect 1750 2785 2800 2800
rect 1750 2765 1765 2785
rect 1785 2765 1815 2785
rect 1835 2765 1865 2785
rect 1885 2765 1915 2785
rect 1935 2765 1965 2785
rect 1985 2765 2015 2785
rect 2035 2765 2065 2785
rect 2085 2765 2115 2785
rect 2135 2765 2165 2785
rect 2185 2765 2215 2785
rect 2235 2765 2265 2785
rect 2285 2765 2315 2785
rect 2335 2765 2365 2785
rect 2385 2765 2415 2785
rect 2435 2765 2465 2785
rect 2485 2765 2515 2785
rect 2535 2765 2565 2785
rect 2585 2765 2615 2785
rect 2635 2765 2665 2785
rect 2685 2765 2715 2785
rect 2735 2765 2765 2785
rect 2785 2765 2800 2785
rect 1750 2750 2800 2765
rect 1750 2735 1800 2750
rect 1750 2715 1765 2735
rect 1785 2715 1800 2735
rect 1750 2685 1800 2715
rect 1750 2665 1765 2685
rect 1785 2665 1800 2685
rect 1750 2635 1800 2665
rect 1750 2615 1765 2635
rect 1785 2615 1800 2635
rect 1750 2585 1800 2615
rect 1750 2565 1765 2585
rect 1785 2565 1800 2585
rect 1750 2535 1800 2565
rect 1750 2515 1765 2535
rect 1785 2515 1800 2535
rect 1750 2485 1800 2515
rect 1750 2465 1765 2485
rect 1785 2465 1800 2485
rect 1750 2435 1800 2465
rect 1750 2415 1765 2435
rect 1785 2415 1800 2435
rect 1750 2385 1800 2415
rect 1750 2365 1765 2385
rect 1785 2365 1800 2385
rect 1750 2335 1800 2365
rect 1750 2315 1765 2335
rect 1785 2315 1800 2335
rect 1750 2285 1800 2315
rect 1750 2265 1765 2285
rect 1785 2265 1800 2285
rect 1750 2235 1800 2265
rect 1750 2215 1765 2235
rect 1785 2215 1800 2235
rect 1750 2185 1800 2215
rect 1750 2165 1765 2185
rect 1785 2165 1800 2185
rect 1750 2135 1800 2165
rect 1750 2115 1765 2135
rect 1785 2115 1800 2135
rect 1750 2085 1800 2115
rect 1750 2065 1765 2085
rect 1785 2065 1800 2085
rect 1750 2035 1800 2065
rect 1750 2015 1765 2035
rect 1785 2015 1800 2035
rect 1750 1985 1800 2015
rect 1850 2685 1900 2700
rect 1850 2665 1865 2685
rect 1885 2665 1900 2685
rect 1850 2635 1900 2665
rect 1850 2615 1865 2635
rect 1885 2615 1900 2635
rect 1850 2585 1900 2615
rect 1850 2565 1865 2585
rect 1885 2565 1900 2585
rect 1850 2535 1900 2565
rect 1850 2515 1865 2535
rect 1885 2515 1900 2535
rect 1850 2485 1900 2515
rect 1850 2465 1865 2485
rect 1885 2465 1900 2485
rect 1850 2435 1900 2465
rect 1850 2415 1865 2435
rect 1885 2415 1900 2435
rect 1850 2385 1900 2415
rect 1850 2365 1865 2385
rect 1885 2365 1900 2385
rect 1850 2335 1900 2365
rect 1850 2315 1865 2335
rect 1885 2315 1900 2335
rect 1850 2285 1900 2315
rect 1850 2265 1865 2285
rect 1885 2265 1900 2285
rect 1850 2235 1900 2265
rect 1850 2215 1865 2235
rect 1885 2215 1900 2235
rect 1850 2185 1900 2215
rect 1850 2165 1865 2185
rect 1885 2165 1900 2185
rect 1850 2135 1900 2165
rect 1850 2115 1865 2135
rect 1885 2115 1900 2135
rect 1850 2085 1900 2115
rect 1850 2065 1865 2085
rect 1885 2065 1900 2085
rect 1850 2035 1900 2065
rect 1850 2015 1865 2035
rect 1885 2015 1900 2035
rect 1850 2000 1900 2015
rect 2050 2685 2100 2700
rect 2050 2665 2065 2685
rect 2085 2665 2100 2685
rect 2050 2635 2100 2665
rect 2050 2615 2065 2635
rect 2085 2615 2100 2635
rect 2050 2585 2100 2615
rect 2050 2565 2065 2585
rect 2085 2565 2100 2585
rect 2050 2535 2100 2565
rect 2050 2515 2065 2535
rect 2085 2515 2100 2535
rect 2050 2485 2100 2515
rect 2050 2465 2065 2485
rect 2085 2465 2100 2485
rect 2050 2435 2100 2465
rect 2050 2415 2065 2435
rect 2085 2415 2100 2435
rect 2050 2385 2100 2415
rect 2050 2365 2065 2385
rect 2085 2365 2100 2385
rect 2050 2335 2100 2365
rect 2050 2315 2065 2335
rect 2085 2315 2100 2335
rect 2050 2285 2100 2315
rect 2050 2265 2065 2285
rect 2085 2265 2100 2285
rect 2050 2235 2100 2265
rect 2050 2215 2065 2235
rect 2085 2215 2100 2235
rect 2050 2185 2100 2215
rect 2050 2165 2065 2185
rect 2085 2165 2100 2185
rect 2050 2135 2100 2165
rect 2050 2115 2065 2135
rect 2085 2115 2100 2135
rect 2050 2085 2100 2115
rect 2050 2065 2065 2085
rect 2085 2065 2100 2085
rect 2050 2035 2100 2065
rect 2050 2015 2065 2035
rect 2085 2015 2100 2035
rect 2050 2000 2100 2015
rect 2250 2685 2300 2750
rect 2750 2735 2800 2750
rect 2750 2715 2765 2735
rect 2785 2715 2800 2735
rect 2250 2665 2265 2685
rect 2285 2665 2300 2685
rect 2250 2635 2300 2665
rect 2250 2615 2265 2635
rect 2285 2615 2300 2635
rect 2250 2585 2300 2615
rect 2250 2565 2265 2585
rect 2285 2565 2300 2585
rect 2250 2535 2300 2565
rect 2250 2515 2265 2535
rect 2285 2515 2300 2535
rect 2250 2485 2300 2515
rect 2250 2465 2265 2485
rect 2285 2465 2300 2485
rect 2250 2435 2300 2465
rect 2250 2415 2265 2435
rect 2285 2415 2300 2435
rect 2250 2385 2300 2415
rect 2250 2365 2265 2385
rect 2285 2365 2300 2385
rect 2250 2335 2300 2365
rect 2250 2315 2265 2335
rect 2285 2315 2300 2335
rect 2250 2285 2300 2315
rect 2250 2265 2265 2285
rect 2285 2265 2300 2285
rect 2250 2235 2300 2265
rect 2250 2215 2265 2235
rect 2285 2215 2300 2235
rect 2250 2185 2300 2215
rect 2250 2165 2265 2185
rect 2285 2165 2300 2185
rect 2250 2135 2300 2165
rect 2250 2115 2265 2135
rect 2285 2115 2300 2135
rect 2250 2085 2300 2115
rect 2250 2065 2265 2085
rect 2285 2065 2300 2085
rect 2250 2035 2300 2065
rect 2250 2015 2265 2035
rect 2285 2015 2300 2035
rect 2250 2000 2300 2015
rect 2450 2685 2500 2700
rect 2450 2665 2465 2685
rect 2485 2665 2500 2685
rect 2450 2635 2500 2665
rect 2450 2615 2465 2635
rect 2485 2615 2500 2635
rect 2450 2585 2500 2615
rect 2450 2565 2465 2585
rect 2485 2565 2500 2585
rect 2450 2535 2500 2565
rect 2450 2515 2465 2535
rect 2485 2515 2500 2535
rect 2450 2485 2500 2515
rect 2450 2465 2465 2485
rect 2485 2465 2500 2485
rect 2450 2435 2500 2465
rect 2450 2415 2465 2435
rect 2485 2415 2500 2435
rect 2450 2385 2500 2415
rect 2450 2365 2465 2385
rect 2485 2365 2500 2385
rect 2450 2335 2500 2365
rect 2450 2315 2465 2335
rect 2485 2315 2500 2335
rect 2450 2285 2500 2315
rect 2450 2265 2465 2285
rect 2485 2265 2500 2285
rect 2450 2235 2500 2265
rect 2450 2215 2465 2235
rect 2485 2215 2500 2235
rect 2450 2185 2500 2215
rect 2450 2165 2465 2185
rect 2485 2165 2500 2185
rect 2450 2135 2500 2165
rect 2450 2115 2465 2135
rect 2485 2115 2500 2135
rect 2450 2085 2500 2115
rect 2450 2065 2465 2085
rect 2485 2065 2500 2085
rect 2450 2035 2500 2065
rect 2450 2015 2465 2035
rect 2485 2015 2500 2035
rect 2450 2000 2500 2015
rect 2650 2685 2700 2700
rect 2650 2665 2665 2685
rect 2685 2665 2700 2685
rect 2650 2635 2700 2665
rect 2650 2615 2665 2635
rect 2685 2615 2700 2635
rect 2650 2585 2700 2615
rect 2650 2565 2665 2585
rect 2685 2565 2700 2585
rect 2650 2535 2700 2565
rect 2650 2515 2665 2535
rect 2685 2515 2700 2535
rect 2650 2485 2700 2515
rect 2650 2465 2665 2485
rect 2685 2465 2700 2485
rect 2650 2435 2700 2465
rect 2650 2415 2665 2435
rect 2685 2415 2700 2435
rect 2650 2385 2700 2415
rect 2650 2365 2665 2385
rect 2685 2365 2700 2385
rect 2650 2335 2700 2365
rect 2650 2315 2665 2335
rect 2685 2315 2700 2335
rect 2650 2285 2700 2315
rect 2650 2265 2665 2285
rect 2685 2265 2700 2285
rect 2650 2235 2700 2265
rect 2650 2215 2665 2235
rect 2685 2215 2700 2235
rect 2650 2185 2700 2215
rect 2650 2165 2665 2185
rect 2685 2165 2700 2185
rect 2650 2135 2700 2165
rect 2650 2115 2665 2135
rect 2685 2115 2700 2135
rect 2650 2085 2700 2115
rect 2650 2065 2665 2085
rect 2685 2065 2700 2085
rect 2650 2035 2700 2065
rect 2650 2015 2665 2035
rect 2685 2015 2700 2035
rect 2650 2000 2700 2015
rect 2750 2685 2800 2715
rect 2750 2665 2765 2685
rect 2785 2665 2800 2685
rect 2750 2635 2800 2665
rect 2750 2615 2765 2635
rect 2785 2615 2800 2635
rect 2750 2585 2800 2615
rect 2750 2565 2765 2585
rect 2785 2565 2800 2585
rect 2750 2535 2800 2565
rect 2750 2515 2765 2535
rect 2785 2515 2800 2535
rect 2750 2485 2800 2515
rect 2750 2465 2765 2485
rect 2785 2465 2800 2485
rect 2750 2435 2800 2465
rect 2750 2415 2765 2435
rect 2785 2415 2800 2435
rect 2750 2385 2800 2415
rect 2750 2365 2765 2385
rect 2785 2365 2800 2385
rect 2750 2335 2800 2365
rect 2750 2315 2765 2335
rect 2785 2315 2800 2335
rect 2750 2285 2800 2315
rect 2750 2265 2765 2285
rect 2785 2265 2800 2285
rect 2750 2235 2800 2265
rect 2750 2215 2765 2235
rect 2785 2215 2800 2235
rect 2750 2185 2800 2215
rect 2750 2165 2765 2185
rect 2785 2165 2800 2185
rect 2750 2135 2800 2165
rect 2750 2115 2765 2135
rect 2785 2115 2800 2135
rect 2750 2085 2800 2115
rect 2750 2065 2765 2085
rect 2785 2065 2800 2085
rect 2750 2035 2800 2065
rect 2750 2015 2765 2035
rect 2785 2015 2800 2035
rect 1750 1965 1765 1985
rect 1785 1965 1800 1985
rect 1750 1935 1800 1965
rect 2750 1985 2800 2015
rect 2750 1965 2765 1985
rect 2785 1965 2800 1985
rect 1750 1915 1765 1935
rect 1785 1915 1800 1935
rect 1750 1885 1800 1915
rect 1900 1935 2050 1950
rect 1900 1915 1915 1935
rect 1935 1915 1965 1935
rect 1985 1915 2015 1935
rect 2035 1915 2050 1935
rect 1900 1900 2050 1915
rect 2100 1935 2250 1950
rect 2100 1915 2115 1935
rect 2135 1915 2165 1935
rect 2185 1915 2215 1935
rect 2235 1915 2250 1935
rect 2100 1900 2250 1915
rect 2300 1935 2450 1950
rect 2300 1915 2315 1935
rect 2335 1915 2365 1935
rect 2385 1915 2415 1935
rect 2435 1915 2450 1935
rect 2300 1900 2450 1915
rect 2500 1935 2650 1950
rect 2500 1915 2515 1935
rect 2535 1915 2565 1935
rect 2585 1915 2615 1935
rect 2635 1915 2650 1935
rect 2500 1900 2650 1915
rect 2750 1935 2800 1965
rect 2750 1915 2765 1935
rect 2785 1915 2800 1935
rect 1750 1865 1765 1885
rect 1785 1865 1800 1885
rect 1750 1835 1800 1865
rect 2750 1885 2800 1915
rect 2750 1865 2765 1885
rect 2785 1865 2800 1885
rect 1750 1815 1765 1835
rect 1785 1815 1800 1835
rect 1750 1785 1800 1815
rect 1750 1765 1765 1785
rect 1785 1765 1800 1785
rect 1750 1735 1800 1765
rect 1750 1715 1765 1735
rect 1785 1715 1800 1735
rect 1750 1685 1800 1715
rect 1750 1665 1765 1685
rect 1785 1665 1800 1685
rect 1750 1635 1800 1665
rect 1750 1615 1765 1635
rect 1785 1615 1800 1635
rect 1750 1585 1800 1615
rect 1750 1565 1765 1585
rect 1785 1565 1800 1585
rect 1750 1535 1800 1565
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1750 1485 1800 1515
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1850 1835 1900 1850
rect 1850 1815 1865 1835
rect 1885 1815 1900 1835
rect 1850 1785 1900 1815
rect 1850 1765 1865 1785
rect 1885 1765 1900 1785
rect 1850 1735 1900 1765
rect 1850 1715 1865 1735
rect 1885 1715 1900 1735
rect 1850 1685 1900 1715
rect 1850 1665 1865 1685
rect 1885 1665 1900 1685
rect 1850 1635 1900 1665
rect 1850 1615 1865 1635
rect 1885 1615 1900 1635
rect 1850 1585 1900 1615
rect 1850 1565 1865 1585
rect 1885 1565 1900 1585
rect 1850 1535 1900 1565
rect 1850 1515 1865 1535
rect 1885 1515 1900 1535
rect 1850 1485 1900 1515
rect 1850 1465 1865 1485
rect 1885 1465 1900 1485
rect 1850 1435 1900 1465
rect 1850 1415 1865 1435
rect 1885 1415 1900 1435
rect 1850 1385 1900 1415
rect 1850 1365 1865 1385
rect 1885 1365 1900 1385
rect 1850 1335 1900 1365
rect 1850 1315 1865 1335
rect 1885 1315 1900 1335
rect 1850 1285 1900 1315
rect 1850 1265 1865 1285
rect 1885 1265 1900 1285
rect 1850 1235 1900 1265
rect 1850 1215 1865 1235
rect 1885 1215 1900 1235
rect 1850 1185 1900 1215
rect 1850 1165 1865 1185
rect 1885 1165 1900 1185
rect 1850 1150 1900 1165
rect 2050 1835 2100 1850
rect 2050 1815 2065 1835
rect 2085 1815 2100 1835
rect 2050 1785 2100 1815
rect 2050 1765 2065 1785
rect 2085 1765 2100 1785
rect 2050 1735 2100 1765
rect 2050 1715 2065 1735
rect 2085 1715 2100 1735
rect 2050 1685 2100 1715
rect 2050 1665 2065 1685
rect 2085 1665 2100 1685
rect 2050 1635 2100 1665
rect 2050 1615 2065 1635
rect 2085 1615 2100 1635
rect 2050 1585 2100 1615
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1150 2100 1165
rect 2250 1835 2300 1850
rect 2250 1815 2265 1835
rect 2285 1815 2300 1835
rect 2250 1785 2300 1815
rect 2250 1765 2265 1785
rect 2285 1765 2300 1785
rect 2250 1735 2300 1765
rect 2250 1715 2265 1735
rect 2285 1715 2300 1735
rect 2250 1685 2300 1715
rect 2250 1665 2265 1685
rect 2285 1665 2300 1685
rect 2250 1635 2300 1665
rect 2250 1615 2265 1635
rect 2285 1615 2300 1635
rect 2250 1585 2300 1615
rect 2250 1565 2265 1585
rect 2285 1565 2300 1585
rect 2250 1535 2300 1565
rect 2250 1515 2265 1535
rect 2285 1515 2300 1535
rect 2250 1485 2300 1515
rect 2250 1465 2265 1485
rect 2285 1465 2300 1485
rect 2250 1435 2300 1465
rect 2250 1415 2265 1435
rect 2285 1415 2300 1435
rect 2250 1385 2300 1415
rect 2250 1365 2265 1385
rect 2285 1365 2300 1385
rect 2250 1335 2300 1365
rect 2250 1315 2265 1335
rect 2285 1315 2300 1335
rect 2250 1285 2300 1315
rect 2250 1265 2265 1285
rect 2285 1265 2300 1285
rect 2250 1235 2300 1265
rect 2250 1215 2265 1235
rect 2285 1215 2300 1235
rect 2250 1185 2300 1215
rect 2250 1165 2265 1185
rect 2285 1165 2300 1185
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1100 1800 1115
rect 2250 1100 2300 1165
rect 2450 1835 2500 1850
rect 2450 1815 2465 1835
rect 2485 1815 2500 1835
rect 2450 1785 2500 1815
rect 2450 1765 2465 1785
rect 2485 1765 2500 1785
rect 2450 1735 2500 1765
rect 2450 1715 2465 1735
rect 2485 1715 2500 1735
rect 2450 1685 2500 1715
rect 2450 1665 2465 1685
rect 2485 1665 2500 1685
rect 2450 1635 2500 1665
rect 2450 1615 2465 1635
rect 2485 1615 2500 1635
rect 2450 1585 2500 1615
rect 2450 1565 2465 1585
rect 2485 1565 2500 1585
rect 2450 1535 2500 1565
rect 2450 1515 2465 1535
rect 2485 1515 2500 1535
rect 2450 1485 2500 1515
rect 2450 1465 2465 1485
rect 2485 1465 2500 1485
rect 2450 1435 2500 1465
rect 2450 1415 2465 1435
rect 2485 1415 2500 1435
rect 2450 1385 2500 1415
rect 2450 1365 2465 1385
rect 2485 1365 2500 1385
rect 2450 1335 2500 1365
rect 2450 1315 2465 1335
rect 2485 1315 2500 1335
rect 2450 1285 2500 1315
rect 2450 1265 2465 1285
rect 2485 1265 2500 1285
rect 2450 1235 2500 1265
rect 2450 1215 2465 1235
rect 2485 1215 2500 1235
rect 2450 1185 2500 1215
rect 2450 1165 2465 1185
rect 2485 1165 2500 1185
rect 2450 1150 2500 1165
rect 2650 1835 2700 1850
rect 2650 1815 2665 1835
rect 2685 1815 2700 1835
rect 2650 1785 2700 1815
rect 2650 1765 2665 1785
rect 2685 1765 2700 1785
rect 2650 1735 2700 1765
rect 2650 1715 2665 1735
rect 2685 1715 2700 1735
rect 2650 1685 2700 1715
rect 2650 1665 2665 1685
rect 2685 1665 2700 1685
rect 2650 1635 2700 1665
rect 2650 1615 2665 1635
rect 2685 1615 2700 1635
rect 2650 1585 2700 1615
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1150 2700 1165
rect 2750 1835 2800 1865
rect 2750 1815 2765 1835
rect 2785 1815 2800 1835
rect 2750 1785 2800 1815
rect 2750 1765 2765 1785
rect 2785 1765 2800 1785
rect 2750 1735 2800 1765
rect 2750 1715 2765 1735
rect 2785 1715 2800 1735
rect 2750 1685 2800 1715
rect 2750 1665 2765 1685
rect 2785 1665 2800 1685
rect 2750 1635 2800 1665
rect 2750 1615 2765 1635
rect 2785 1615 2800 1635
rect 2750 1585 2800 1615
rect 2750 1565 2765 1585
rect 2785 1565 2800 1585
rect 2750 1535 2800 1565
rect 2750 1515 2765 1535
rect 2785 1515 2800 1535
rect 2750 1485 2800 1515
rect 2750 1465 2765 1485
rect 2785 1465 2800 1485
rect 2750 1435 2800 1465
rect 2750 1415 2765 1435
rect 2785 1415 2800 1435
rect 2750 1385 2800 1415
rect 2750 1365 2765 1385
rect 2785 1365 2800 1385
rect 2750 1335 2800 1365
rect 2750 1315 2765 1335
rect 2785 1315 2800 1335
rect 2750 1285 2800 1315
rect 2750 1265 2765 1285
rect 2785 1265 2800 1285
rect 2750 1235 2800 1265
rect 2750 1215 2765 1235
rect 2785 1215 2800 1235
rect 2750 1185 2800 1215
rect 2750 1165 2765 1185
rect 2785 1165 2800 1185
rect 2750 1135 2800 1165
rect 2750 1115 2765 1135
rect 2785 1115 2800 1135
rect 2750 1100 2800 1115
rect 1750 1085 2800 1100
rect 1750 1065 1765 1085
rect 1785 1065 1815 1085
rect 1835 1065 1865 1085
rect 1885 1065 1915 1085
rect 1935 1065 1965 1085
rect 1985 1065 2015 1085
rect 2035 1065 2065 1085
rect 2085 1065 2115 1085
rect 2135 1065 2165 1085
rect 2185 1065 2215 1085
rect 2235 1065 2265 1085
rect 2285 1065 2315 1085
rect 2335 1065 2365 1085
rect 2385 1065 2415 1085
rect 2435 1065 2465 1085
rect 2485 1065 2515 1085
rect 2535 1065 2565 1085
rect 2585 1065 2615 1085
rect 2635 1065 2665 1085
rect 2685 1065 2715 1085
rect 2735 1065 2765 1085
rect 2785 1065 2800 1085
rect 1750 1050 2800 1065
rect 2900 2785 2950 2815
rect 2900 2765 2915 2785
rect 2935 2765 2950 2785
rect 2900 2735 2950 2765
rect 2900 2715 2915 2735
rect 2935 2715 2950 2735
rect 2900 2685 2950 2715
rect 2900 2665 2915 2685
rect 2935 2665 2950 2685
rect 2900 2635 2950 2665
rect 2900 2615 2915 2635
rect 2935 2615 2950 2635
rect 2900 2585 2950 2615
rect 2900 2565 2915 2585
rect 2935 2565 2950 2585
rect 2900 2535 2950 2565
rect 2900 2515 2915 2535
rect 2935 2515 2950 2535
rect 2900 2485 2950 2515
rect 2900 2465 2915 2485
rect 2935 2465 2950 2485
rect 2900 2435 2950 2465
rect 2900 2415 2915 2435
rect 2935 2415 2950 2435
rect 2900 2385 2950 2415
rect 2900 2365 2915 2385
rect 2935 2365 2950 2385
rect 2900 2335 2950 2365
rect 2900 2315 2915 2335
rect 2935 2315 2950 2335
rect 2900 2285 2950 2315
rect 2900 2265 2915 2285
rect 2935 2265 2950 2285
rect 2900 2235 2950 2265
rect 2900 2215 2915 2235
rect 2935 2215 2950 2235
rect 2900 2185 2950 2215
rect 2900 2165 2915 2185
rect 2935 2165 2950 2185
rect 2900 2135 2950 2165
rect 2900 2115 2915 2135
rect 2935 2115 2950 2135
rect 2900 2085 2950 2115
rect 2900 2065 2915 2085
rect 2935 2065 2950 2085
rect 2900 2035 2950 2065
rect 2900 2015 2915 2035
rect 2935 2015 2950 2035
rect 2900 1985 2950 2015
rect 2900 1965 2915 1985
rect 2935 1965 2950 1985
rect 2900 1935 2950 1965
rect 2900 1915 2915 1935
rect 2935 1915 2950 1935
rect 2900 1885 2950 1915
rect 2900 1865 2915 1885
rect 2935 1865 2950 1885
rect 2900 1835 2950 1865
rect 2900 1815 2915 1835
rect 2935 1815 2950 1835
rect 2900 1785 2950 1815
rect 2900 1765 2915 1785
rect 2935 1765 2950 1785
rect 2900 1735 2950 1765
rect 2900 1715 2915 1735
rect 2935 1715 2950 1735
rect 2900 1685 2950 1715
rect 2900 1665 2915 1685
rect 2935 1665 2950 1685
rect 2900 1635 2950 1665
rect 2900 1615 2915 1635
rect 2935 1615 2950 1635
rect 2900 1585 2950 1615
rect 2900 1565 2915 1585
rect 2935 1565 2950 1585
rect 2900 1535 2950 1565
rect 2900 1515 2915 1535
rect 2935 1515 2950 1535
rect 2900 1485 2950 1515
rect 2900 1465 2915 1485
rect 2935 1465 2950 1485
rect 2900 1435 2950 1465
rect 2900 1415 2915 1435
rect 2935 1415 2950 1435
rect 2900 1385 2950 1415
rect 2900 1365 2915 1385
rect 2935 1365 2950 1385
rect 2900 1335 2950 1365
rect 2900 1315 2915 1335
rect 2935 1315 2950 1335
rect 2900 1285 2950 1315
rect 2900 1265 2915 1285
rect 2935 1265 2950 1285
rect 2900 1235 2950 1265
rect 2900 1215 2915 1235
rect 2935 1215 2950 1235
rect 2900 1185 2950 1215
rect 2900 1165 2915 1185
rect 2935 1165 2950 1185
rect 2900 1135 2950 1165
rect 2900 1115 2915 1135
rect 2935 1115 2950 1135
rect 2900 1085 2950 1115
rect 2900 1065 2915 1085
rect 2935 1065 2950 1085
rect 1600 1015 1615 1035
rect 1635 1015 1650 1035
rect 1600 985 1650 1015
rect 1600 965 1615 985
rect 1635 965 1650 985
rect 1600 950 1650 965
rect 2900 1035 2950 1065
rect 2900 1015 2915 1035
rect 2935 1015 2950 1035
rect 2900 985 2950 1015
rect 2900 965 2915 985
rect 2935 965 2950 985
rect 2900 950 2950 965
rect 1600 935 2950 950
rect 1600 915 1615 935
rect 1635 915 1665 935
rect 1685 915 1715 935
rect 1735 915 1765 935
rect 1785 915 1815 935
rect 1835 915 1865 935
rect 1885 915 1915 935
rect 1935 915 1965 935
rect 1985 915 2015 935
rect 2035 915 2065 935
rect 2085 915 2115 935
rect 2135 915 2165 935
rect 2185 915 2215 935
rect 2235 915 2265 935
rect 2285 915 2315 935
rect 2335 915 2365 935
rect 2385 915 2415 935
rect 2435 915 2465 935
rect 2485 915 2515 935
rect 2535 915 2565 935
rect 2585 915 2615 935
rect 2635 915 2665 935
rect 2685 915 2715 935
rect 2735 915 2765 935
rect 2785 915 2815 935
rect 2835 915 2865 935
rect 2885 915 2915 935
rect 2935 915 2950 935
rect 1600 900 2950 915
rect 1600 885 1650 900
rect 1600 865 1615 885
rect 1635 865 1650 885
rect 1600 835 1650 865
rect 2900 885 2950 900
rect 2900 865 2915 885
rect 2935 865 2950 885
rect 1600 815 1615 835
rect 1635 815 1650 835
rect 1600 785 1650 815
rect 1900 835 2050 850
rect 1900 815 1915 835
rect 1935 815 1965 835
rect 1985 815 2015 835
rect 2035 815 2050 835
rect 1900 800 2050 815
rect 2100 835 2250 850
rect 2100 815 2115 835
rect 2135 815 2165 835
rect 2185 815 2215 835
rect 2235 815 2250 835
rect 2100 800 2250 815
rect 2300 835 2450 850
rect 2300 815 2315 835
rect 2335 815 2365 835
rect 2385 815 2415 835
rect 2435 815 2450 835
rect 2300 800 2450 815
rect 2500 835 2650 850
rect 2500 815 2515 835
rect 2535 815 2565 835
rect 2585 815 2615 835
rect 2635 815 2650 835
rect 2500 800 2650 815
rect 2900 835 2950 865
rect 2900 815 2915 835
rect 2935 815 2950 835
rect 1600 765 1615 785
rect 1635 765 1650 785
rect 1600 735 1650 765
rect 2900 785 2950 815
rect 2900 765 2915 785
rect 2935 765 2950 785
rect 1600 715 1615 735
rect 1635 715 1650 735
rect 1600 685 1650 715
rect 1600 665 1615 685
rect 1635 665 1650 685
rect 1600 635 1650 665
rect 1600 615 1615 635
rect 1635 615 1650 635
rect 1600 585 1650 615
rect 1600 565 1615 585
rect 1635 565 1650 585
rect 1600 535 1650 565
rect 1600 515 1615 535
rect 1635 515 1650 535
rect 1600 485 1650 515
rect 1600 465 1615 485
rect 1635 465 1650 485
rect 1600 435 1650 465
rect 1600 415 1615 435
rect 1635 415 1650 435
rect 1600 385 1650 415
rect 1600 365 1615 385
rect 1635 365 1650 385
rect 1600 335 1650 365
rect 1600 315 1615 335
rect 1635 315 1650 335
rect 1600 285 1650 315
rect 1600 265 1615 285
rect 1635 265 1650 285
rect 1600 235 1650 265
rect 1850 735 1900 750
rect 1850 715 1865 735
rect 1885 715 1900 735
rect 1850 685 1900 715
rect 1850 665 1865 685
rect 1885 665 1900 685
rect 1850 635 1900 665
rect 1850 615 1865 635
rect 1885 615 1900 635
rect 1850 585 1900 615
rect 1850 565 1865 585
rect 1885 565 1900 585
rect 1850 535 1900 565
rect 1850 515 1865 535
rect 1885 515 1900 535
rect 1850 485 1900 515
rect 1850 465 1865 485
rect 1885 465 1900 485
rect 1850 435 1900 465
rect 1850 415 1865 435
rect 1885 415 1900 435
rect 1850 385 1900 415
rect 1850 365 1865 385
rect 1885 365 1900 385
rect 1850 335 1900 365
rect 1850 315 1865 335
rect 1885 315 1900 335
rect 1850 285 1900 315
rect 1850 265 1865 285
rect 1885 265 1900 285
rect 1850 250 1900 265
rect 1950 735 2000 750
rect 1950 715 1965 735
rect 1985 715 2000 735
rect 1950 685 2000 715
rect 1950 665 1965 685
rect 1985 665 2000 685
rect 1950 635 2000 665
rect 1950 615 1965 635
rect 1985 615 2000 635
rect 1950 585 2000 615
rect 1950 565 1965 585
rect 1985 565 2000 585
rect 1950 535 2000 565
rect 1950 515 1965 535
rect 1985 515 2000 535
rect 1950 485 2000 515
rect 1950 465 1965 485
rect 1985 465 2000 485
rect 1950 435 2000 465
rect 1950 415 1965 435
rect 1985 415 2000 435
rect 1950 385 2000 415
rect 1950 365 1965 385
rect 1985 365 2000 385
rect 1950 335 2000 365
rect 1950 315 1965 335
rect 1985 315 2000 335
rect 1950 285 2000 315
rect 1950 265 1965 285
rect 1985 265 2000 285
rect 1950 250 2000 265
rect 2050 735 2100 750
rect 2050 715 2065 735
rect 2085 715 2100 735
rect 2050 685 2100 715
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 2050 635 2100 665
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 250 2100 265
rect 2150 735 2200 750
rect 2150 715 2165 735
rect 2185 715 2200 735
rect 2150 685 2200 715
rect 2150 665 2165 685
rect 2185 665 2200 685
rect 2150 635 2200 665
rect 2150 615 2165 635
rect 2185 615 2200 635
rect 2150 585 2200 615
rect 2150 565 2165 585
rect 2185 565 2200 585
rect 2150 535 2200 565
rect 2150 515 2165 535
rect 2185 515 2200 535
rect 2150 485 2200 515
rect 2150 465 2165 485
rect 2185 465 2200 485
rect 2150 435 2200 465
rect 2150 415 2165 435
rect 2185 415 2200 435
rect 2150 385 2200 415
rect 2150 365 2165 385
rect 2185 365 2200 385
rect 2150 335 2200 365
rect 2150 315 2165 335
rect 2185 315 2200 335
rect 2150 285 2200 315
rect 2150 265 2165 285
rect 2185 265 2200 285
rect 2150 250 2200 265
rect 2250 735 2300 750
rect 2250 715 2265 735
rect 2285 715 2300 735
rect 2250 685 2300 715
rect 2250 665 2265 685
rect 2285 665 2300 685
rect 2250 635 2300 665
rect 2250 615 2265 635
rect 2285 615 2300 635
rect 2250 585 2300 615
rect 2250 565 2265 585
rect 2285 565 2300 585
rect 2250 535 2300 565
rect 2250 515 2265 535
rect 2285 515 2300 535
rect 2250 485 2300 515
rect 2250 465 2265 485
rect 2285 465 2300 485
rect 2250 435 2300 465
rect 2250 415 2265 435
rect 2285 415 2300 435
rect 2250 385 2300 415
rect 2250 365 2265 385
rect 2285 365 2300 385
rect 2250 335 2300 365
rect 2250 315 2265 335
rect 2285 315 2300 335
rect 2250 285 2300 315
rect 2250 265 2265 285
rect 2285 265 2300 285
rect 1600 215 1615 235
rect 1635 215 1650 235
rect 1600 200 1650 215
rect 2250 200 2300 265
rect 2350 735 2400 750
rect 2350 715 2365 735
rect 2385 715 2400 735
rect 2350 685 2400 715
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 250 2400 265
rect 2450 735 2500 750
rect 2450 715 2465 735
rect 2485 715 2500 735
rect 2450 685 2500 715
rect 2450 665 2465 685
rect 2485 665 2500 685
rect 2450 635 2500 665
rect 2450 615 2465 635
rect 2485 615 2500 635
rect 2450 585 2500 615
rect 2450 565 2465 585
rect 2485 565 2500 585
rect 2450 535 2500 565
rect 2450 515 2465 535
rect 2485 515 2500 535
rect 2450 485 2500 515
rect 2450 465 2465 485
rect 2485 465 2500 485
rect 2450 435 2500 465
rect 2450 415 2465 435
rect 2485 415 2500 435
rect 2450 385 2500 415
rect 2450 365 2465 385
rect 2485 365 2500 385
rect 2450 335 2500 365
rect 2450 315 2465 335
rect 2485 315 2500 335
rect 2450 285 2500 315
rect 2450 265 2465 285
rect 2485 265 2500 285
rect 2450 250 2500 265
rect 2550 735 2600 750
rect 2550 715 2565 735
rect 2585 715 2600 735
rect 2550 685 2600 715
rect 2550 665 2565 685
rect 2585 665 2600 685
rect 2550 635 2600 665
rect 2550 615 2565 635
rect 2585 615 2600 635
rect 2550 585 2600 615
rect 2550 565 2565 585
rect 2585 565 2600 585
rect 2550 535 2600 565
rect 2550 515 2565 535
rect 2585 515 2600 535
rect 2550 485 2600 515
rect 2550 465 2565 485
rect 2585 465 2600 485
rect 2550 435 2600 465
rect 2550 415 2565 435
rect 2585 415 2600 435
rect 2550 385 2600 415
rect 2550 365 2565 385
rect 2585 365 2600 385
rect 2550 335 2600 365
rect 2550 315 2565 335
rect 2585 315 2600 335
rect 2550 285 2600 315
rect 2550 265 2565 285
rect 2585 265 2600 285
rect 2550 250 2600 265
rect 2650 735 2700 750
rect 2650 715 2665 735
rect 2685 715 2700 735
rect 2650 685 2700 715
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 635 2700 665
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 250 2700 265
rect 2900 735 2950 765
rect 2900 715 2915 735
rect 2935 715 2950 735
rect 2900 685 2950 715
rect 2900 665 2915 685
rect 2935 665 2950 685
rect 2900 635 2950 665
rect 2900 615 2915 635
rect 2935 615 2950 635
rect 2900 585 2950 615
rect 2900 565 2915 585
rect 2935 565 2950 585
rect 2900 535 2950 565
rect 2900 515 2915 535
rect 2935 515 2950 535
rect 2900 485 2950 515
rect 2900 465 2915 485
rect 2935 465 2950 485
rect 2900 435 2950 465
rect 2900 415 2915 435
rect 2935 415 2950 435
rect 2900 385 2950 415
rect 2900 365 2915 385
rect 2935 365 2950 385
rect 2900 335 2950 365
rect 2900 315 2915 335
rect 2935 315 2950 335
rect 2900 285 2950 315
rect 2900 265 2915 285
rect 2935 265 2950 285
rect 2900 235 2950 265
rect 2900 215 2915 235
rect 2935 215 2950 235
rect 2900 200 2950 215
rect 1600 185 2950 200
rect 1600 165 1615 185
rect 1635 165 1665 185
rect 1685 165 1715 185
rect 1735 165 1765 185
rect 1785 165 1815 185
rect 1835 165 1865 185
rect 1885 165 1915 185
rect 1935 165 1965 185
rect 1985 165 2015 185
rect 2035 165 2065 185
rect 2085 165 2115 185
rect 2135 165 2165 185
rect 2185 165 2215 185
rect 2235 165 2265 185
rect 2285 165 2315 185
rect 2335 165 2365 185
rect 2385 165 2415 185
rect 2435 165 2465 185
rect 2485 165 2515 185
rect 2535 165 2565 185
rect 2585 165 2615 185
rect 2635 165 2665 185
rect 2685 165 2715 185
rect 2735 165 2765 185
rect 2785 165 2815 185
rect 2835 165 2865 185
rect 2885 165 2915 185
rect 2935 165 2950 185
rect 1600 150 2950 165
rect 3050 3685 3100 3715
rect 3050 3665 3065 3685
rect 3085 3665 3100 3685
rect 3050 3635 3100 3665
rect 3050 3615 3065 3635
rect 3085 3615 3100 3635
rect 3050 3585 3100 3615
rect 3050 3565 3065 3585
rect 3085 3565 3100 3585
rect 3050 3535 3100 3565
rect 3050 3515 3065 3535
rect 3085 3515 3100 3535
rect 3050 3485 3100 3515
rect 3050 3465 3065 3485
rect 3085 3465 3100 3485
rect 3050 3435 3100 3465
rect 3050 3415 3065 3435
rect 3085 3415 3100 3435
rect 3050 3385 3100 3415
rect 3050 3365 3065 3385
rect 3085 3365 3100 3385
rect 3050 3335 3100 3365
rect 3050 3315 3065 3335
rect 3085 3315 3100 3335
rect 3050 3285 3100 3315
rect 3050 3265 3065 3285
rect 3085 3265 3100 3285
rect 3050 3235 3100 3265
rect 3050 3215 3065 3235
rect 3085 3215 3100 3235
rect 3050 3185 3100 3215
rect 3050 3165 3065 3185
rect 3085 3165 3100 3185
rect 3050 3135 3100 3165
rect 3050 3115 3065 3135
rect 3085 3115 3100 3135
rect 3050 3085 3100 3115
rect 3050 3065 3065 3085
rect 3085 3065 3100 3085
rect 3050 3035 3100 3065
rect 3050 3015 3065 3035
rect 3085 3015 3100 3035
rect 3050 2985 3100 3015
rect 3050 2965 3065 2985
rect 3085 2965 3100 2985
rect 3050 2935 3100 2965
rect 3050 2915 3065 2935
rect 3085 2915 3100 2935
rect 3050 2885 3100 2915
rect 3050 2865 3065 2885
rect 3085 2865 3100 2885
rect 3050 2835 3100 2865
rect 3050 2815 3065 2835
rect 3085 2815 3100 2835
rect 3050 2785 3100 2815
rect 3050 2765 3065 2785
rect 3085 2765 3100 2785
rect 3050 2735 3100 2765
rect 3050 2715 3065 2735
rect 3085 2715 3100 2735
rect 3050 2685 3100 2715
rect 3050 2665 3065 2685
rect 3085 2665 3100 2685
rect 3050 2635 3100 2665
rect 3050 2615 3065 2635
rect 3085 2615 3100 2635
rect 3050 2585 3100 2615
rect 3050 2565 3065 2585
rect 3085 2565 3100 2585
rect 3050 2535 3100 2565
rect 3050 2515 3065 2535
rect 3085 2515 3100 2535
rect 3050 2485 3100 2515
rect 3050 2465 3065 2485
rect 3085 2465 3100 2485
rect 3050 2435 3100 2465
rect 3050 2415 3065 2435
rect 3085 2415 3100 2435
rect 3050 2385 3100 2415
rect 3050 2365 3065 2385
rect 3085 2365 3100 2385
rect 3050 2335 3100 2365
rect 3050 2315 3065 2335
rect 3085 2315 3100 2335
rect 3050 2285 3100 2315
rect 3050 2265 3065 2285
rect 3085 2265 3100 2285
rect 3050 2235 3100 2265
rect 3050 2215 3065 2235
rect 3085 2215 3100 2235
rect 3050 2185 3100 2215
rect 3050 2165 3065 2185
rect 3085 2165 3100 2185
rect 3050 2135 3100 2165
rect 3050 2115 3065 2135
rect 3085 2115 3100 2135
rect 3050 2085 3100 2115
rect 3050 2065 3065 2085
rect 3085 2065 3100 2085
rect 3050 2035 3100 2065
rect 3050 2015 3065 2035
rect 3085 2015 3100 2035
rect 3050 1985 3100 2015
rect 3050 1965 3065 1985
rect 3085 1965 3100 1985
rect 3050 1935 3100 1965
rect 3050 1915 3065 1935
rect 3085 1915 3100 1935
rect 3050 1885 3100 1915
rect 3050 1865 3065 1885
rect 3085 1865 3100 1885
rect 3050 1835 3100 1865
rect 3050 1815 3065 1835
rect 3085 1815 3100 1835
rect 3050 1785 3100 1815
rect 3050 1765 3065 1785
rect 3085 1765 3100 1785
rect 3050 1735 3100 1765
rect 3050 1715 3065 1735
rect 3085 1715 3100 1735
rect 3050 1685 3100 1715
rect 3050 1665 3065 1685
rect 3085 1665 3100 1685
rect 3050 1635 3100 1665
rect 3050 1615 3065 1635
rect 3085 1615 3100 1635
rect 3050 1585 3100 1615
rect 3050 1565 3065 1585
rect 3085 1565 3100 1585
rect 3050 1535 3100 1565
rect 3050 1515 3065 1535
rect 3085 1515 3100 1535
rect 3050 1485 3100 1515
rect 3050 1465 3065 1485
rect 3085 1465 3100 1485
rect 3050 1435 3100 1465
rect 3050 1415 3065 1435
rect 3085 1415 3100 1435
rect 3050 1385 3100 1415
rect 3050 1365 3065 1385
rect 3085 1365 3100 1385
rect 3050 1335 3100 1365
rect 3050 1315 3065 1335
rect 3085 1315 3100 1335
rect 3050 1285 3100 1315
rect 3050 1265 3065 1285
rect 3085 1265 3100 1285
rect 3050 1235 3100 1265
rect 3050 1215 3065 1235
rect 3085 1215 3100 1235
rect 3050 1185 3100 1215
rect 3050 1165 3065 1185
rect 3085 1165 3100 1185
rect 3050 1135 3100 1165
rect 3050 1115 3065 1135
rect 3085 1115 3100 1135
rect 3050 1085 3100 1115
rect 3050 1065 3065 1085
rect 3085 1065 3100 1085
rect 3050 1035 3100 1065
rect 3050 1015 3065 1035
rect 3085 1015 3100 1035
rect 3050 985 3100 1015
rect 3050 965 3065 985
rect 3085 965 3100 985
rect 3050 935 3100 965
rect 3050 915 3065 935
rect 3085 915 3100 935
rect 3050 885 3100 915
rect 3050 865 3065 885
rect 3085 865 3100 885
rect 3050 835 3100 865
rect 3050 815 3065 835
rect 3085 815 3100 835
rect 3050 785 3100 815
rect 3050 765 3065 785
rect 3085 765 3100 785
rect 3050 735 3100 765
rect 3050 715 3065 735
rect 3085 715 3100 735
rect 3050 685 3100 715
rect 3050 665 3065 685
rect 3085 665 3100 685
rect 3050 635 3100 665
rect 3050 615 3065 635
rect 3085 615 3100 635
rect 3050 585 3100 615
rect 3050 565 3065 585
rect 3085 565 3100 585
rect 3050 535 3100 565
rect 3050 515 3065 535
rect 3085 515 3100 535
rect 3050 485 3100 515
rect 3050 465 3065 485
rect 3085 465 3100 485
rect 3050 435 3100 465
rect 3050 415 3065 435
rect 3085 415 3100 435
rect 3050 385 3100 415
rect 3050 365 3065 385
rect 3085 365 3100 385
rect 3050 335 3100 365
rect 3050 315 3065 335
rect 3085 315 3100 335
rect 3050 285 3100 315
rect 3050 265 3065 285
rect 3085 265 3100 285
rect 3050 235 3100 265
rect 3050 215 3065 235
rect 3085 215 3100 235
rect 3050 185 3100 215
rect 3050 165 3065 185
rect 3085 165 3100 185
rect 1450 115 1465 135
rect 1485 115 1500 135
rect 1450 85 1500 115
rect 1450 65 1465 85
rect 1485 65 1500 85
rect 1450 50 1500 65
rect 3050 135 3100 165
rect 3050 115 3065 135
rect 3085 115 3100 135
rect 3050 85 3100 115
rect 3050 65 3065 85
rect 3085 65 3100 85
rect 3050 50 3100 65
rect 1450 35 3100 50
rect 1450 15 1465 35
rect 1485 15 1515 35
rect 1535 15 1565 35
rect 1585 15 1615 35
rect 1635 15 1665 35
rect 1685 15 1715 35
rect 1735 15 1765 35
rect 1785 15 1815 35
rect 1835 15 1865 35
rect 1885 15 1915 35
rect 1935 15 1965 35
rect 1985 15 2015 35
rect 2035 15 2065 35
rect 2085 15 2115 35
rect 2135 15 2165 35
rect 2185 15 2215 35
rect 2235 15 2265 35
rect 2285 15 2315 35
rect 2335 15 2365 35
rect 2385 15 2415 35
rect 2435 15 2465 35
rect 2485 15 2515 35
rect 2535 15 2565 35
rect 2585 15 2615 35
rect 2635 15 2665 35
rect 2685 15 2715 35
rect 2735 15 2765 35
rect 2785 15 2815 35
rect 2835 15 2865 35
rect 2885 15 2915 35
rect 2935 15 2965 35
rect 2985 15 3015 35
rect 3035 15 3065 35
rect 3085 15 3100 35
rect 1450 0 3100 15
<< viali >>
rect 1865 3565 1885 3585
rect 1865 3515 1885 3535
rect 1865 3465 1885 3485
rect 1865 3415 1885 3435
rect 1865 3365 1885 3385
rect 1865 3315 1885 3335
rect 1865 3265 1885 3285
rect 1865 3215 1885 3235
rect 1865 3165 1885 3185
rect 1865 3115 1885 3135
rect 1965 3565 1985 3585
rect 1965 3515 1985 3535
rect 1965 3465 1985 3485
rect 1965 3415 1985 3435
rect 1965 3365 1985 3385
rect 1965 3315 1985 3335
rect 1965 3265 1985 3285
rect 1965 3215 1985 3235
rect 1965 3165 1985 3185
rect 1965 3115 1985 3135
rect 2065 3565 2085 3585
rect 2065 3515 2085 3535
rect 2065 3465 2085 3485
rect 2065 3415 2085 3435
rect 2065 3365 2085 3385
rect 2065 3315 2085 3335
rect 2065 3265 2085 3285
rect 2065 3215 2085 3235
rect 2165 3565 2185 3585
rect 2165 3515 2185 3535
rect 2165 3465 2185 3485
rect 2165 3415 2185 3435
rect 2165 3365 2185 3385
rect 2165 3315 2185 3335
rect 2165 3265 2185 3285
rect 2165 3215 2185 3235
rect 2165 3165 2185 3185
rect 2165 3115 2185 3135
rect 2365 3565 2385 3585
rect 2365 3515 2385 3535
rect 2365 3465 2385 3485
rect 2365 3415 2385 3435
rect 2365 3365 2385 3385
rect 2365 3315 2385 3335
rect 2365 3265 2385 3285
rect 2365 3215 2385 3235
rect 2365 3165 2385 3185
rect 2365 3115 2385 3135
rect 2465 3565 2485 3585
rect 2465 3515 2485 3535
rect 2465 3465 2485 3485
rect 2465 3415 2485 3435
rect 2465 3365 2485 3385
rect 2465 3315 2485 3335
rect 2465 3265 2485 3285
rect 2465 3215 2485 3235
rect 2565 3565 2585 3585
rect 2565 3515 2585 3535
rect 2565 3465 2585 3485
rect 2565 3415 2585 3435
rect 2565 3365 2585 3385
rect 2565 3315 2585 3335
rect 2565 3265 2585 3285
rect 2565 3215 2585 3235
rect 2565 3165 2585 3185
rect 2565 3115 2585 3135
rect 2665 3565 2685 3585
rect 2665 3515 2685 3535
rect 2665 3465 2685 3485
rect 2665 3415 2685 3435
rect 2665 3365 2685 3385
rect 2665 3315 2685 3335
rect 2665 3265 2685 3285
rect 2665 3215 2685 3235
rect 2665 3165 2685 3185
rect 2665 3115 2685 3135
rect 1965 3015 1985 3035
rect 2165 3015 2185 3035
rect 2365 3015 2385 3035
rect 2565 3015 2585 3035
rect 1865 2665 1885 2685
rect 1865 2615 1885 2635
rect 1865 2565 1885 2585
rect 1865 2515 1885 2535
rect 1865 2465 1885 2485
rect 1865 2415 1885 2435
rect 1865 2365 1885 2385
rect 1865 2315 1885 2335
rect 1865 2265 1885 2285
rect 1865 2215 1885 2235
rect 1865 2165 1885 2185
rect 1865 2115 1885 2135
rect 1865 2065 1885 2085
rect 1865 2015 1885 2035
rect 2065 2665 2085 2685
rect 2065 2615 2085 2635
rect 2065 2565 2085 2585
rect 2065 2515 2085 2535
rect 2065 2465 2085 2485
rect 2065 2415 2085 2435
rect 2065 2365 2085 2385
rect 2065 2315 2085 2335
rect 2065 2265 2085 2285
rect 2065 2215 2085 2235
rect 2065 2165 2085 2185
rect 2065 2115 2085 2135
rect 2065 2065 2085 2085
rect 2065 2015 2085 2035
rect 2465 2665 2485 2685
rect 2465 2615 2485 2635
rect 2465 2565 2485 2585
rect 2465 2515 2485 2535
rect 2465 2465 2485 2485
rect 2465 2415 2485 2435
rect 2465 2365 2485 2385
rect 2465 2315 2485 2335
rect 2465 2265 2485 2285
rect 2465 2215 2485 2235
rect 2465 2165 2485 2185
rect 2465 2115 2485 2135
rect 2465 2065 2485 2085
rect 2465 2015 2485 2035
rect 2665 2665 2685 2685
rect 2665 2615 2685 2635
rect 2665 2565 2685 2585
rect 2665 2515 2685 2535
rect 2665 2465 2685 2485
rect 2665 2415 2685 2435
rect 2665 2365 2685 2385
rect 2665 2315 2685 2335
rect 2665 2265 2685 2285
rect 2665 2215 2685 2235
rect 2665 2165 2685 2185
rect 2665 2115 2685 2135
rect 2665 2065 2685 2085
rect 2665 2015 2685 2035
rect 1965 1915 1985 1935
rect 2165 1915 2185 1935
rect 2365 1915 2385 1935
rect 2565 1915 2585 1935
rect 1865 1815 1885 1835
rect 1865 1765 1885 1785
rect 1865 1715 1885 1735
rect 1865 1665 1885 1685
rect 1865 1615 1885 1635
rect 1865 1565 1885 1585
rect 1865 1515 1885 1535
rect 1865 1465 1885 1485
rect 1865 1415 1885 1435
rect 1865 1365 1885 1385
rect 1865 1315 1885 1335
rect 1865 1265 1885 1285
rect 1865 1215 1885 1235
rect 1865 1165 1885 1185
rect 2065 1815 2085 1835
rect 2065 1765 2085 1785
rect 2065 1715 2085 1735
rect 2065 1665 2085 1685
rect 2065 1615 2085 1635
rect 2065 1565 2085 1585
rect 2065 1515 2085 1535
rect 2065 1465 2085 1485
rect 2065 1415 2085 1435
rect 2065 1365 2085 1385
rect 2065 1315 2085 1335
rect 2065 1265 2085 1285
rect 2065 1215 2085 1235
rect 2065 1165 2085 1185
rect 2465 1815 2485 1835
rect 2465 1765 2485 1785
rect 2465 1715 2485 1735
rect 2465 1665 2485 1685
rect 2465 1615 2485 1635
rect 2465 1565 2485 1585
rect 2465 1515 2485 1535
rect 2465 1465 2485 1485
rect 2465 1415 2485 1435
rect 2465 1365 2485 1385
rect 2465 1315 2485 1335
rect 2465 1265 2485 1285
rect 2465 1215 2485 1235
rect 2465 1165 2485 1185
rect 2665 1815 2685 1835
rect 2665 1765 2685 1785
rect 2665 1715 2685 1735
rect 2665 1665 2685 1685
rect 2665 1615 2685 1635
rect 2665 1565 2685 1585
rect 2665 1515 2685 1535
rect 2665 1465 2685 1485
rect 2665 1415 2685 1435
rect 2665 1365 2685 1385
rect 2665 1315 2685 1335
rect 2665 1265 2685 1285
rect 2665 1215 2685 1235
rect 2665 1165 2685 1185
rect 1965 815 1985 835
rect 2165 815 2185 835
rect 2365 815 2385 835
rect 2565 815 2585 835
rect 1865 715 1885 735
rect 1865 665 1885 685
rect 1865 615 1885 635
rect 1865 565 1885 585
rect 1865 515 1885 535
rect 1865 465 1885 485
rect 1865 415 1885 435
rect 1865 365 1885 385
rect 1865 315 1885 335
rect 1865 265 1885 285
rect 1965 715 1985 735
rect 1965 665 1985 685
rect 1965 615 1985 635
rect 1965 565 1985 585
rect 1965 515 1985 535
rect 1965 465 1985 485
rect 1965 415 1985 435
rect 1965 365 1985 385
rect 1965 315 1985 335
rect 1965 265 1985 285
rect 2065 615 2085 635
rect 2065 565 2085 585
rect 2065 515 2085 535
rect 2065 465 2085 485
rect 2065 415 2085 435
rect 2065 365 2085 385
rect 2065 315 2085 335
rect 2065 265 2085 285
rect 2165 715 2185 735
rect 2165 665 2185 685
rect 2165 615 2185 635
rect 2165 565 2185 585
rect 2165 515 2185 535
rect 2165 465 2185 485
rect 2165 415 2185 435
rect 2165 365 2185 385
rect 2165 315 2185 335
rect 2165 265 2185 285
rect 2365 715 2385 735
rect 2365 665 2385 685
rect 2365 615 2385 635
rect 2365 565 2385 585
rect 2365 515 2385 535
rect 2365 465 2385 485
rect 2365 415 2385 435
rect 2365 365 2385 385
rect 2365 315 2385 335
rect 2365 265 2385 285
rect 2465 615 2485 635
rect 2465 565 2485 585
rect 2465 515 2485 535
rect 2465 465 2485 485
rect 2465 415 2485 435
rect 2465 365 2485 385
rect 2465 315 2485 335
rect 2465 265 2485 285
rect 2565 715 2585 735
rect 2565 665 2585 685
rect 2565 615 2585 635
rect 2565 565 2585 585
rect 2565 515 2585 535
rect 2565 465 2585 485
rect 2565 415 2585 435
rect 2565 365 2585 385
rect 2565 315 2585 335
rect 2565 265 2585 285
rect 2665 715 2685 735
rect 2665 665 2685 685
rect 2665 615 2685 635
rect 2665 565 2685 585
rect 2665 515 2685 535
rect 2665 465 2685 485
rect 2665 415 2685 435
rect 2665 365 2685 385
rect 2665 315 2685 335
rect 2665 265 2685 285
<< metal1 >>
rect 1850 3740 1900 3750
rect 1850 3710 1860 3740
rect 1890 3710 1900 3740
rect 1850 3640 1900 3710
rect 1850 3610 1860 3640
rect 1890 3610 1900 3640
rect 1850 3585 1900 3610
rect 2050 3740 2100 3750
rect 2050 3710 2060 3740
rect 2090 3710 2100 3740
rect 2050 3640 2100 3710
rect 2050 3610 2060 3640
rect 2090 3610 2100 3640
rect 1850 3565 1865 3585
rect 1885 3565 1900 3585
rect 1850 3540 1900 3565
rect 1850 3510 1860 3540
rect 1890 3510 1900 3540
rect 1850 3485 1900 3510
rect 1850 3465 1865 3485
rect 1885 3465 1900 3485
rect 1850 3440 1900 3465
rect 1850 3410 1860 3440
rect 1890 3410 1900 3440
rect 1850 3385 1900 3410
rect 1850 3365 1865 3385
rect 1885 3365 1900 3385
rect 1850 3340 1900 3365
rect 1850 3310 1860 3340
rect 1890 3310 1900 3340
rect 1850 3285 1900 3310
rect 1850 3265 1865 3285
rect 1885 3265 1900 3285
rect 1850 3240 1900 3265
rect 1850 3210 1860 3240
rect 1890 3210 1900 3240
rect 1850 3185 1900 3210
rect 1850 3165 1865 3185
rect 1885 3165 1900 3185
rect 1850 3140 1900 3165
rect 1850 3110 1860 3140
rect 1890 3110 1900 3140
rect 1850 3100 1900 3110
rect 1950 3585 2000 3600
rect 1950 3565 1965 3585
rect 1985 3565 2000 3585
rect 1950 3535 2000 3565
rect 1950 3515 1965 3535
rect 1985 3515 2000 3535
rect 1950 3485 2000 3515
rect 1950 3465 1965 3485
rect 1985 3465 2000 3485
rect 1950 3435 2000 3465
rect 1950 3415 1965 3435
rect 1985 3415 2000 3435
rect 1950 3385 2000 3415
rect 1950 3365 1965 3385
rect 1985 3365 2000 3385
rect 1950 3335 2000 3365
rect 1950 3315 1965 3335
rect 1985 3315 2000 3335
rect 1950 3285 2000 3315
rect 1950 3265 1965 3285
rect 1985 3265 2000 3285
rect 1950 3235 2000 3265
rect 1950 3215 1965 3235
rect 1985 3215 2000 3235
rect 1950 3185 2000 3215
rect 2050 3585 2100 3610
rect 2450 3740 2500 3750
rect 2450 3710 2460 3740
rect 2490 3710 2500 3740
rect 2450 3640 2500 3710
rect 2450 3610 2460 3640
rect 2490 3610 2500 3640
rect 2050 3565 2065 3585
rect 2085 3565 2100 3585
rect 2050 3540 2100 3565
rect 2050 3510 2060 3540
rect 2090 3510 2100 3540
rect 2050 3485 2100 3510
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3440 2100 3465
rect 2050 3410 2060 3440
rect 2090 3410 2100 3440
rect 2050 3385 2100 3410
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3340 2100 3365
rect 2050 3310 2060 3340
rect 2090 3310 2100 3340
rect 2050 3285 2100 3310
rect 2050 3265 2065 3285
rect 2085 3265 2100 3285
rect 2050 3240 2100 3265
rect 2050 3210 2060 3240
rect 2090 3210 2100 3240
rect 2050 3200 2100 3210
rect 2150 3585 2200 3600
rect 2150 3565 2165 3585
rect 2185 3565 2200 3585
rect 2150 3535 2200 3565
rect 2150 3515 2165 3535
rect 2185 3515 2200 3535
rect 2150 3485 2200 3515
rect 2150 3465 2165 3485
rect 2185 3465 2200 3485
rect 2150 3435 2200 3465
rect 2150 3415 2165 3435
rect 2185 3415 2200 3435
rect 2150 3385 2200 3415
rect 2150 3365 2165 3385
rect 2185 3365 2200 3385
rect 2150 3335 2200 3365
rect 2150 3315 2165 3335
rect 2185 3315 2200 3335
rect 2150 3285 2200 3315
rect 2150 3265 2165 3285
rect 2185 3265 2200 3285
rect 2150 3235 2200 3265
rect 2150 3215 2165 3235
rect 2185 3215 2200 3235
rect 1950 3165 1965 3185
rect 1985 3165 2000 3185
rect 1950 3150 2000 3165
rect 2150 3185 2200 3215
rect 2150 3165 2165 3185
rect 2185 3165 2200 3185
rect 2150 3150 2200 3165
rect 1950 3135 2200 3150
rect 1950 3115 1965 3135
rect 1985 3115 2165 3135
rect 2185 3115 2200 3135
rect 1950 3100 2200 3115
rect 2350 3585 2400 3600
rect 2350 3565 2365 3585
rect 2385 3565 2400 3585
rect 2350 3535 2400 3565
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3285 2400 3315
rect 2350 3265 2365 3285
rect 2385 3265 2400 3285
rect 2350 3235 2400 3265
rect 2350 3215 2365 3235
rect 2385 3215 2400 3235
rect 2350 3185 2400 3215
rect 2450 3585 2500 3610
rect 2650 3740 2700 3750
rect 2650 3710 2660 3740
rect 2690 3710 2700 3740
rect 2650 3640 2700 3710
rect 2650 3610 2660 3640
rect 2690 3610 2700 3640
rect 2450 3565 2465 3585
rect 2485 3565 2500 3585
rect 2450 3540 2500 3565
rect 2450 3510 2460 3540
rect 2490 3510 2500 3540
rect 2450 3485 2500 3510
rect 2450 3465 2465 3485
rect 2485 3465 2500 3485
rect 2450 3440 2500 3465
rect 2450 3410 2460 3440
rect 2490 3410 2500 3440
rect 2450 3385 2500 3410
rect 2450 3365 2465 3385
rect 2485 3365 2500 3385
rect 2450 3340 2500 3365
rect 2450 3310 2460 3340
rect 2490 3310 2500 3340
rect 2450 3285 2500 3310
rect 2450 3265 2465 3285
rect 2485 3265 2500 3285
rect 2450 3240 2500 3265
rect 2450 3210 2460 3240
rect 2490 3210 2500 3240
rect 2450 3200 2500 3210
rect 2550 3585 2600 3600
rect 2550 3565 2565 3585
rect 2585 3565 2600 3585
rect 2550 3535 2600 3565
rect 2550 3515 2565 3535
rect 2585 3515 2600 3535
rect 2550 3485 2600 3515
rect 2550 3465 2565 3485
rect 2585 3465 2600 3485
rect 2550 3435 2600 3465
rect 2550 3415 2565 3435
rect 2585 3415 2600 3435
rect 2550 3385 2600 3415
rect 2550 3365 2565 3385
rect 2585 3365 2600 3385
rect 2550 3335 2600 3365
rect 2550 3315 2565 3335
rect 2585 3315 2600 3335
rect 2550 3285 2600 3315
rect 2550 3265 2565 3285
rect 2585 3265 2600 3285
rect 2550 3235 2600 3265
rect 2550 3215 2565 3235
rect 2585 3215 2600 3235
rect 2350 3165 2365 3185
rect 2385 3165 2400 3185
rect 2350 3150 2400 3165
rect 2550 3185 2600 3215
rect 2550 3165 2565 3185
rect 2585 3165 2600 3185
rect 2550 3150 2600 3165
rect 2350 3135 2600 3150
rect 2350 3115 2365 3135
rect 2385 3115 2565 3135
rect 2585 3115 2600 3135
rect 2350 3100 2600 3115
rect 2650 3585 2700 3610
rect 2650 3565 2665 3585
rect 2685 3565 2700 3585
rect 2650 3540 2700 3565
rect 2650 3510 2660 3540
rect 2690 3510 2700 3540
rect 2650 3485 2700 3510
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3440 2700 3465
rect 2650 3410 2660 3440
rect 2690 3410 2700 3440
rect 2650 3385 2700 3410
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3340 2700 3365
rect 2650 3310 2660 3340
rect 2690 3310 2700 3340
rect 2650 3285 2700 3310
rect 2650 3265 2665 3285
rect 2685 3265 2700 3285
rect 2650 3240 2700 3265
rect 2650 3210 2660 3240
rect 2690 3210 2700 3240
rect 2650 3185 2700 3210
rect 2650 3165 2665 3185
rect 2685 3165 2700 3185
rect 2650 3140 2700 3165
rect 2650 3110 2660 3140
rect 2690 3110 2700 3140
rect 2650 3100 2700 3110
rect 1950 3040 2000 3050
rect 1950 3010 1960 3040
rect 1990 3010 2000 3040
rect 1950 3000 2000 3010
rect 1850 2840 1900 2850
rect 1850 2810 1860 2840
rect 1890 2810 1900 2840
rect 1850 2685 1900 2810
rect 1850 2665 1865 2685
rect 1885 2665 1900 2685
rect 1850 2635 1900 2665
rect 1850 2615 1865 2635
rect 1885 2615 1900 2635
rect 1850 2585 1900 2615
rect 1850 2565 1865 2585
rect 1885 2565 1900 2585
rect 1850 2535 1900 2565
rect 1850 2515 1865 2535
rect 1885 2515 1900 2535
rect 1850 2485 1900 2515
rect 1850 2465 1865 2485
rect 1885 2465 1900 2485
rect 1850 2440 1900 2465
rect 1850 2410 1860 2440
rect 1890 2410 1900 2440
rect 1850 2385 1900 2410
rect 1850 2365 1865 2385
rect 1885 2365 1900 2385
rect 1850 2335 1900 2365
rect 1850 2315 1865 2335
rect 1885 2315 1900 2335
rect 1850 2285 1900 2315
rect 1850 2265 1865 2285
rect 1885 2265 1900 2285
rect 1850 2240 1900 2265
rect 1850 2210 1860 2240
rect 1890 2210 1900 2240
rect 1850 2185 1900 2210
rect 1850 2165 1865 2185
rect 1885 2165 1900 2185
rect 1850 2135 1900 2165
rect 1850 2115 1865 2135
rect 1885 2115 1900 2135
rect 1850 2085 1900 2115
rect 1850 2065 1865 2085
rect 1885 2065 1900 2085
rect 1850 2040 1900 2065
rect 1850 2010 1860 2040
rect 1890 2010 1900 2040
rect 1850 1840 1900 2010
rect 2050 2685 2100 3100
rect 2150 3040 2200 3050
rect 2150 3010 2160 3040
rect 2190 3010 2200 3040
rect 2150 3000 2200 3010
rect 2350 3040 2400 3050
rect 2350 3010 2360 3040
rect 2390 3010 2400 3040
rect 2350 3000 2400 3010
rect 2050 2665 2065 2685
rect 2085 2665 2100 2685
rect 2050 2635 2100 2665
rect 2050 2615 2065 2635
rect 2085 2615 2100 2635
rect 2050 2585 2100 2615
rect 2050 2565 2065 2585
rect 2085 2565 2100 2585
rect 2050 2535 2100 2565
rect 2050 2515 2065 2535
rect 2085 2515 2100 2535
rect 2050 2485 2100 2515
rect 2050 2465 2065 2485
rect 2085 2465 2100 2485
rect 2050 2435 2100 2465
rect 2050 2415 2065 2435
rect 2085 2415 2100 2435
rect 2050 2385 2100 2415
rect 2050 2365 2065 2385
rect 2085 2365 2100 2385
rect 2050 2335 2100 2365
rect 2050 2315 2065 2335
rect 2085 2315 2100 2335
rect 2050 2285 2100 2315
rect 2050 2265 2065 2285
rect 2085 2265 2100 2285
rect 2050 2235 2100 2265
rect 2050 2215 2065 2235
rect 2085 2215 2100 2235
rect 2050 2185 2100 2215
rect 2050 2165 2065 2185
rect 2085 2165 2100 2185
rect 2050 2135 2100 2165
rect 2050 2115 2065 2135
rect 2085 2115 2100 2135
rect 2050 2085 2100 2115
rect 2050 2065 2065 2085
rect 2085 2065 2100 2085
rect 2050 2035 2100 2065
rect 2050 2015 2065 2035
rect 2085 2015 2100 2035
rect 2050 1950 2100 2015
rect 2450 2685 2500 3100
rect 2550 3040 2600 3050
rect 2550 3010 2560 3040
rect 2590 3010 2600 3040
rect 2550 3000 2600 3010
rect 2450 2665 2465 2685
rect 2485 2665 2500 2685
rect 2450 2635 2500 2665
rect 2450 2615 2465 2635
rect 2485 2615 2500 2635
rect 2450 2585 2500 2615
rect 2450 2565 2465 2585
rect 2485 2565 2500 2585
rect 2450 2535 2500 2565
rect 2450 2515 2465 2535
rect 2485 2515 2500 2535
rect 2450 2485 2500 2515
rect 2450 2465 2465 2485
rect 2485 2465 2500 2485
rect 2450 2435 2500 2465
rect 2450 2415 2465 2435
rect 2485 2415 2500 2435
rect 2450 2385 2500 2415
rect 2450 2365 2465 2385
rect 2485 2365 2500 2385
rect 2450 2335 2500 2365
rect 2450 2315 2465 2335
rect 2485 2315 2500 2335
rect 2450 2285 2500 2315
rect 2450 2265 2465 2285
rect 2485 2265 2500 2285
rect 2450 2235 2500 2265
rect 2450 2215 2465 2235
rect 2485 2215 2500 2235
rect 2450 2185 2500 2215
rect 2450 2165 2465 2185
rect 2485 2165 2500 2185
rect 2450 2135 2500 2165
rect 2450 2115 2465 2135
rect 2485 2115 2500 2135
rect 2450 2085 2500 2115
rect 2450 2065 2465 2085
rect 2485 2065 2500 2085
rect 2450 2035 2500 2065
rect 2450 2015 2465 2035
rect 2485 2015 2500 2035
rect 2450 1950 2500 2015
rect 2650 2840 2700 2850
rect 2650 2810 2660 2840
rect 2690 2810 2700 2840
rect 2650 2685 2700 2810
rect 2650 2665 2665 2685
rect 2685 2665 2700 2685
rect 2650 2635 2700 2665
rect 2650 2615 2665 2635
rect 2685 2615 2700 2635
rect 2650 2585 2700 2615
rect 2650 2565 2665 2585
rect 2685 2565 2700 2585
rect 2650 2535 2700 2565
rect 2650 2515 2665 2535
rect 2685 2515 2700 2535
rect 2650 2485 2700 2515
rect 2650 2465 2665 2485
rect 2685 2465 2700 2485
rect 2650 2440 2700 2465
rect 2650 2410 2660 2440
rect 2690 2410 2700 2440
rect 2650 2385 2700 2410
rect 2650 2365 2665 2385
rect 2685 2365 2700 2385
rect 2650 2335 2700 2365
rect 2650 2315 2665 2335
rect 2685 2315 2700 2335
rect 2650 2285 2700 2315
rect 2650 2265 2665 2285
rect 2685 2265 2700 2285
rect 2650 2240 2700 2265
rect 2650 2210 2660 2240
rect 2690 2210 2700 2240
rect 2650 2185 2700 2210
rect 2650 2165 2665 2185
rect 2685 2165 2700 2185
rect 2650 2135 2700 2165
rect 2650 2115 2665 2135
rect 2685 2115 2700 2135
rect 2650 2085 2700 2115
rect 2650 2065 2665 2085
rect 2685 2065 2700 2085
rect 2650 2040 2700 2065
rect 2650 2010 2660 2040
rect 2690 2010 2700 2040
rect 1950 1940 2000 1950
rect 1950 1910 1960 1940
rect 1990 1910 2000 1940
rect 1950 1900 2000 1910
rect 2050 1940 2500 1950
rect 2050 1910 2160 1940
rect 2190 1910 2360 1940
rect 2390 1910 2500 1940
rect 2050 1900 2500 1910
rect 2550 1940 2600 1950
rect 2550 1910 2560 1940
rect 2590 1910 2600 1940
rect 2550 1900 2600 1910
rect 1850 1810 1860 1840
rect 1890 1810 1900 1840
rect 1850 1785 1900 1810
rect 1850 1765 1865 1785
rect 1885 1765 1900 1785
rect 1850 1735 1900 1765
rect 1850 1715 1865 1735
rect 1885 1715 1900 1735
rect 1850 1685 1900 1715
rect 1850 1665 1865 1685
rect 1885 1665 1900 1685
rect 1850 1640 1900 1665
rect 1850 1610 1860 1640
rect 1890 1610 1900 1640
rect 1850 1585 1900 1610
rect 1850 1565 1865 1585
rect 1885 1565 1900 1585
rect 1850 1535 1900 1565
rect 1850 1515 1865 1535
rect 1885 1515 1900 1535
rect 1850 1485 1900 1515
rect 1850 1465 1865 1485
rect 1885 1465 1900 1485
rect 1850 1440 1900 1465
rect 1850 1410 1860 1440
rect 1890 1410 1900 1440
rect 1850 1385 1900 1410
rect 1850 1365 1865 1385
rect 1885 1365 1900 1385
rect 1850 1335 1900 1365
rect 1850 1315 1865 1335
rect 1885 1315 1900 1335
rect 1850 1285 1900 1315
rect 1850 1265 1865 1285
rect 1885 1265 1900 1285
rect 1850 1235 1900 1265
rect 1850 1215 1865 1235
rect 1885 1215 1900 1235
rect 1850 1185 1900 1215
rect 1850 1165 1865 1185
rect 1885 1165 1900 1185
rect 1850 1040 1900 1165
rect 1850 1010 1860 1040
rect 1890 1010 1900 1040
rect 1850 1000 1900 1010
rect 2050 1835 2100 1900
rect 2050 1815 2065 1835
rect 2085 1815 2100 1835
rect 2050 1785 2100 1815
rect 2050 1765 2065 1785
rect 2085 1765 2100 1785
rect 2050 1735 2100 1765
rect 2050 1715 2065 1735
rect 2085 1715 2100 1735
rect 2050 1685 2100 1715
rect 2050 1665 2065 1685
rect 2085 1665 2100 1685
rect 2050 1635 2100 1665
rect 2050 1615 2065 1635
rect 2085 1615 2100 1635
rect 2050 1585 2100 1615
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 1950 840 2000 850
rect 1950 810 1960 840
rect 1990 810 2000 840
rect 1950 800 2000 810
rect 2050 750 2100 1165
rect 2450 1835 2500 1900
rect 2450 1815 2465 1835
rect 2485 1815 2500 1835
rect 2450 1785 2500 1815
rect 2450 1765 2465 1785
rect 2485 1765 2500 1785
rect 2450 1735 2500 1765
rect 2450 1715 2465 1735
rect 2485 1715 2500 1735
rect 2450 1685 2500 1715
rect 2450 1665 2465 1685
rect 2485 1665 2500 1685
rect 2450 1635 2500 1665
rect 2450 1615 2465 1635
rect 2485 1615 2500 1635
rect 2450 1585 2500 1615
rect 2450 1565 2465 1585
rect 2485 1565 2500 1585
rect 2450 1535 2500 1565
rect 2450 1515 2465 1535
rect 2485 1515 2500 1535
rect 2450 1485 2500 1515
rect 2450 1465 2465 1485
rect 2485 1465 2500 1485
rect 2450 1435 2500 1465
rect 2450 1415 2465 1435
rect 2485 1415 2500 1435
rect 2450 1385 2500 1415
rect 2450 1365 2465 1385
rect 2485 1365 2500 1385
rect 2450 1335 2500 1365
rect 2450 1315 2465 1335
rect 2485 1315 2500 1335
rect 2450 1285 2500 1315
rect 2450 1265 2465 1285
rect 2485 1265 2500 1285
rect 2450 1235 2500 1265
rect 2450 1215 2465 1235
rect 2485 1215 2500 1235
rect 2450 1185 2500 1215
rect 2450 1165 2465 1185
rect 2485 1165 2500 1185
rect 2150 840 2200 850
rect 2150 810 2160 840
rect 2190 810 2200 840
rect 2150 800 2200 810
rect 2350 840 2400 850
rect 2350 810 2360 840
rect 2390 810 2400 840
rect 2350 800 2400 810
rect 2450 750 2500 1165
rect 2650 1840 2700 2010
rect 2650 1810 2660 1840
rect 2690 1810 2700 1840
rect 2650 1785 2700 1810
rect 2650 1765 2665 1785
rect 2685 1765 2700 1785
rect 2650 1735 2700 1765
rect 2650 1715 2665 1735
rect 2685 1715 2700 1735
rect 2650 1685 2700 1715
rect 2650 1665 2665 1685
rect 2685 1665 2700 1685
rect 2650 1640 2700 1665
rect 2650 1610 2660 1640
rect 2690 1610 2700 1640
rect 2650 1585 2700 1610
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1440 2700 1465
rect 2650 1410 2660 1440
rect 2690 1410 2700 1440
rect 2650 1385 2700 1410
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1040 2700 1165
rect 2650 1010 2660 1040
rect 2690 1010 2700 1040
rect 2650 1000 2700 1010
rect 2550 840 2600 850
rect 2550 810 2560 840
rect 2590 810 2600 840
rect 2550 800 2600 810
rect 1850 740 1900 750
rect 1850 710 1860 740
rect 1890 710 1900 740
rect 1850 685 1900 710
rect 1850 665 1865 685
rect 1885 665 1900 685
rect 1850 640 1900 665
rect 1850 610 1860 640
rect 1890 610 1900 640
rect 1850 585 1900 610
rect 1850 565 1865 585
rect 1885 565 1900 585
rect 1850 540 1900 565
rect 1850 510 1860 540
rect 1890 510 1900 540
rect 1850 485 1900 510
rect 1850 465 1865 485
rect 1885 465 1900 485
rect 1850 440 1900 465
rect 1850 410 1860 440
rect 1890 410 1900 440
rect 1850 385 1900 410
rect 1850 365 1865 385
rect 1885 365 1900 385
rect 1850 340 1900 365
rect 1850 310 1860 340
rect 1890 310 1900 340
rect 1850 285 1900 310
rect 1850 265 1865 285
rect 1885 265 1900 285
rect 1850 240 1900 265
rect 1950 735 2200 750
rect 1950 715 1965 735
rect 1985 715 2165 735
rect 2185 715 2200 735
rect 1950 700 2200 715
rect 1950 685 2000 700
rect 1950 665 1965 685
rect 1985 665 2000 685
rect 1950 635 2000 665
rect 2150 685 2200 700
rect 2150 665 2165 685
rect 2185 665 2200 685
rect 1950 615 1965 635
rect 1985 615 2000 635
rect 1950 585 2000 615
rect 1950 565 1965 585
rect 1985 565 2000 585
rect 1950 535 2000 565
rect 1950 515 1965 535
rect 1985 515 2000 535
rect 1950 485 2000 515
rect 1950 465 1965 485
rect 1985 465 2000 485
rect 1950 435 2000 465
rect 1950 415 1965 435
rect 1985 415 2000 435
rect 1950 385 2000 415
rect 1950 365 1965 385
rect 1985 365 2000 385
rect 1950 335 2000 365
rect 1950 315 1965 335
rect 1985 315 2000 335
rect 1950 285 2000 315
rect 1950 265 1965 285
rect 1985 265 2000 285
rect 1950 250 2000 265
rect 2050 640 2100 650
rect 2050 610 2060 640
rect 2090 610 2100 640
rect 2050 585 2100 610
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 540 2100 565
rect 2050 510 2060 540
rect 2090 510 2100 540
rect 2050 485 2100 510
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 440 2100 465
rect 2050 410 2060 440
rect 2090 410 2100 440
rect 2050 385 2100 410
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 340 2100 365
rect 2050 310 2060 340
rect 2090 310 2100 340
rect 2050 285 2100 310
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 1850 210 1860 240
rect 1890 210 1900 240
rect 1850 140 1900 210
rect 1850 110 1860 140
rect 1890 110 1900 140
rect 1850 100 1900 110
rect 2050 240 2100 265
rect 2150 635 2200 665
rect 2150 615 2165 635
rect 2185 615 2200 635
rect 2150 585 2200 615
rect 2150 565 2165 585
rect 2185 565 2200 585
rect 2150 535 2200 565
rect 2150 515 2165 535
rect 2185 515 2200 535
rect 2150 485 2200 515
rect 2150 465 2165 485
rect 2185 465 2200 485
rect 2150 435 2200 465
rect 2150 415 2165 435
rect 2185 415 2200 435
rect 2150 385 2200 415
rect 2150 365 2165 385
rect 2185 365 2200 385
rect 2150 335 2200 365
rect 2150 315 2165 335
rect 2185 315 2200 335
rect 2150 285 2200 315
rect 2150 265 2165 285
rect 2185 265 2200 285
rect 2150 250 2200 265
rect 2350 735 2600 750
rect 2350 715 2365 735
rect 2385 715 2565 735
rect 2585 715 2600 735
rect 2350 700 2600 715
rect 2350 685 2400 700
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2550 685 2600 700
rect 2550 665 2565 685
rect 2585 665 2600 685
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 250 2400 265
rect 2450 640 2500 650
rect 2450 610 2460 640
rect 2490 610 2500 640
rect 2450 585 2500 610
rect 2450 565 2465 585
rect 2485 565 2500 585
rect 2450 540 2500 565
rect 2450 510 2460 540
rect 2490 510 2500 540
rect 2450 485 2500 510
rect 2450 465 2465 485
rect 2485 465 2500 485
rect 2450 440 2500 465
rect 2450 410 2460 440
rect 2490 410 2500 440
rect 2450 385 2500 410
rect 2450 365 2465 385
rect 2485 365 2500 385
rect 2450 340 2500 365
rect 2450 310 2460 340
rect 2490 310 2500 340
rect 2450 285 2500 310
rect 2450 265 2465 285
rect 2485 265 2500 285
rect 2050 210 2060 240
rect 2090 210 2100 240
rect 2050 140 2100 210
rect 2050 110 2060 140
rect 2090 110 2100 140
rect 2050 100 2100 110
rect 2450 240 2500 265
rect 2550 635 2600 665
rect 2550 615 2565 635
rect 2585 615 2600 635
rect 2550 585 2600 615
rect 2550 565 2565 585
rect 2585 565 2600 585
rect 2550 535 2600 565
rect 2550 515 2565 535
rect 2585 515 2600 535
rect 2550 485 2600 515
rect 2550 465 2565 485
rect 2585 465 2600 485
rect 2550 435 2600 465
rect 2550 415 2565 435
rect 2585 415 2600 435
rect 2550 385 2600 415
rect 2550 365 2565 385
rect 2585 365 2600 385
rect 2550 335 2600 365
rect 2550 315 2565 335
rect 2585 315 2600 335
rect 2550 285 2600 315
rect 2550 265 2565 285
rect 2585 265 2600 285
rect 2550 250 2600 265
rect 2650 740 2700 750
rect 2650 710 2660 740
rect 2690 710 2700 740
rect 2650 685 2700 710
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 640 2700 665
rect 2650 610 2660 640
rect 2690 610 2700 640
rect 2650 585 2700 610
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 540 2700 565
rect 2650 510 2660 540
rect 2690 510 2700 540
rect 2650 485 2700 510
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 440 2700 465
rect 2650 410 2660 440
rect 2690 410 2700 440
rect 2650 385 2700 410
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 340 2700 365
rect 2650 310 2660 340
rect 2690 310 2700 340
rect 2650 285 2700 310
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2450 210 2460 240
rect 2490 210 2500 240
rect 2450 140 2500 210
rect 2450 110 2460 140
rect 2490 110 2500 140
rect 2450 100 2500 110
rect 2650 240 2700 265
rect 2650 210 2660 240
rect 2690 210 2700 240
rect 2650 140 2700 210
rect 2650 110 2660 140
rect 2690 110 2700 140
rect 2650 100 2700 110
<< via1 >>
rect 1860 3710 1890 3740
rect 1860 3610 1890 3640
rect 2060 3710 2090 3740
rect 2060 3610 2090 3640
rect 1860 3535 1890 3540
rect 1860 3515 1865 3535
rect 1865 3515 1885 3535
rect 1885 3515 1890 3535
rect 1860 3510 1890 3515
rect 1860 3435 1890 3440
rect 1860 3415 1865 3435
rect 1865 3415 1885 3435
rect 1885 3415 1890 3435
rect 1860 3410 1890 3415
rect 1860 3335 1890 3340
rect 1860 3315 1865 3335
rect 1865 3315 1885 3335
rect 1885 3315 1890 3335
rect 1860 3310 1890 3315
rect 1860 3235 1890 3240
rect 1860 3215 1865 3235
rect 1865 3215 1885 3235
rect 1885 3215 1890 3235
rect 1860 3210 1890 3215
rect 1860 3135 1890 3140
rect 1860 3115 1865 3135
rect 1865 3115 1885 3135
rect 1885 3115 1890 3135
rect 1860 3110 1890 3115
rect 2460 3710 2490 3740
rect 2460 3610 2490 3640
rect 2060 3535 2090 3540
rect 2060 3515 2065 3535
rect 2065 3515 2085 3535
rect 2085 3515 2090 3535
rect 2060 3510 2090 3515
rect 2060 3435 2090 3440
rect 2060 3415 2065 3435
rect 2065 3415 2085 3435
rect 2085 3415 2090 3435
rect 2060 3410 2090 3415
rect 2060 3335 2090 3340
rect 2060 3315 2065 3335
rect 2065 3315 2085 3335
rect 2085 3315 2090 3335
rect 2060 3310 2090 3315
rect 2060 3235 2090 3240
rect 2060 3215 2065 3235
rect 2065 3215 2085 3235
rect 2085 3215 2090 3235
rect 2060 3210 2090 3215
rect 2660 3710 2690 3740
rect 2660 3610 2690 3640
rect 2460 3535 2490 3540
rect 2460 3515 2465 3535
rect 2465 3515 2485 3535
rect 2485 3515 2490 3535
rect 2460 3510 2490 3515
rect 2460 3435 2490 3440
rect 2460 3415 2465 3435
rect 2465 3415 2485 3435
rect 2485 3415 2490 3435
rect 2460 3410 2490 3415
rect 2460 3335 2490 3340
rect 2460 3315 2465 3335
rect 2465 3315 2485 3335
rect 2485 3315 2490 3335
rect 2460 3310 2490 3315
rect 2460 3235 2490 3240
rect 2460 3215 2465 3235
rect 2465 3215 2485 3235
rect 2485 3215 2490 3235
rect 2460 3210 2490 3215
rect 2660 3535 2690 3540
rect 2660 3515 2665 3535
rect 2665 3515 2685 3535
rect 2685 3515 2690 3535
rect 2660 3510 2690 3515
rect 2660 3435 2690 3440
rect 2660 3415 2665 3435
rect 2665 3415 2685 3435
rect 2685 3415 2690 3435
rect 2660 3410 2690 3415
rect 2660 3335 2690 3340
rect 2660 3315 2665 3335
rect 2665 3315 2685 3335
rect 2685 3315 2690 3335
rect 2660 3310 2690 3315
rect 2660 3235 2690 3240
rect 2660 3215 2665 3235
rect 2665 3215 2685 3235
rect 2685 3215 2690 3235
rect 2660 3210 2690 3215
rect 2660 3135 2690 3140
rect 2660 3115 2665 3135
rect 2665 3115 2685 3135
rect 2685 3115 2690 3135
rect 2660 3110 2690 3115
rect 1960 3035 1990 3040
rect 1960 3015 1965 3035
rect 1965 3015 1985 3035
rect 1985 3015 1990 3035
rect 1960 3010 1990 3015
rect 1860 2810 1890 2840
rect 1860 2435 1890 2440
rect 1860 2415 1865 2435
rect 1865 2415 1885 2435
rect 1885 2415 1890 2435
rect 1860 2410 1890 2415
rect 1860 2235 1890 2240
rect 1860 2215 1865 2235
rect 1865 2215 1885 2235
rect 1885 2215 1890 2235
rect 1860 2210 1890 2215
rect 1860 2035 1890 2040
rect 1860 2015 1865 2035
rect 1865 2015 1885 2035
rect 1885 2015 1890 2035
rect 1860 2010 1890 2015
rect 2160 3035 2190 3040
rect 2160 3015 2165 3035
rect 2165 3015 2185 3035
rect 2185 3015 2190 3035
rect 2160 3010 2190 3015
rect 2360 3035 2390 3040
rect 2360 3015 2365 3035
rect 2365 3015 2385 3035
rect 2385 3015 2390 3035
rect 2360 3010 2390 3015
rect 2560 3035 2590 3040
rect 2560 3015 2565 3035
rect 2565 3015 2585 3035
rect 2585 3015 2590 3035
rect 2560 3010 2590 3015
rect 2660 2810 2690 2840
rect 2660 2435 2690 2440
rect 2660 2415 2665 2435
rect 2665 2415 2685 2435
rect 2685 2415 2690 2435
rect 2660 2410 2690 2415
rect 2660 2235 2690 2240
rect 2660 2215 2665 2235
rect 2665 2215 2685 2235
rect 2685 2215 2690 2235
rect 2660 2210 2690 2215
rect 2660 2035 2690 2040
rect 2660 2015 2665 2035
rect 2665 2015 2685 2035
rect 2685 2015 2690 2035
rect 2660 2010 2690 2015
rect 1960 1935 1990 1940
rect 1960 1915 1965 1935
rect 1965 1915 1985 1935
rect 1985 1915 1990 1935
rect 1960 1910 1990 1915
rect 2160 1935 2190 1940
rect 2160 1915 2165 1935
rect 2165 1915 2185 1935
rect 2185 1915 2190 1935
rect 2160 1910 2190 1915
rect 2360 1935 2390 1940
rect 2360 1915 2365 1935
rect 2365 1915 2385 1935
rect 2385 1915 2390 1935
rect 2360 1910 2390 1915
rect 2560 1935 2590 1940
rect 2560 1915 2565 1935
rect 2565 1915 2585 1935
rect 2585 1915 2590 1935
rect 2560 1910 2590 1915
rect 1860 1835 1890 1840
rect 1860 1815 1865 1835
rect 1865 1815 1885 1835
rect 1885 1815 1890 1835
rect 1860 1810 1890 1815
rect 1860 1635 1890 1640
rect 1860 1615 1865 1635
rect 1865 1615 1885 1635
rect 1885 1615 1890 1635
rect 1860 1610 1890 1615
rect 1860 1435 1890 1440
rect 1860 1415 1865 1435
rect 1865 1415 1885 1435
rect 1885 1415 1890 1435
rect 1860 1410 1890 1415
rect 1860 1010 1890 1040
rect 1960 835 1990 840
rect 1960 815 1965 835
rect 1965 815 1985 835
rect 1985 815 1990 835
rect 1960 810 1990 815
rect 2160 835 2190 840
rect 2160 815 2165 835
rect 2165 815 2185 835
rect 2185 815 2190 835
rect 2160 810 2190 815
rect 2360 835 2390 840
rect 2360 815 2365 835
rect 2365 815 2385 835
rect 2385 815 2390 835
rect 2360 810 2390 815
rect 2660 1835 2690 1840
rect 2660 1815 2665 1835
rect 2665 1815 2685 1835
rect 2685 1815 2690 1835
rect 2660 1810 2690 1815
rect 2660 1635 2690 1640
rect 2660 1615 2665 1635
rect 2665 1615 2685 1635
rect 2685 1615 2690 1635
rect 2660 1610 2690 1615
rect 2660 1435 2690 1440
rect 2660 1415 2665 1435
rect 2665 1415 2685 1435
rect 2685 1415 2690 1435
rect 2660 1410 2690 1415
rect 2660 1010 2690 1040
rect 2560 835 2590 840
rect 2560 815 2565 835
rect 2565 815 2585 835
rect 2585 815 2590 835
rect 2560 810 2590 815
rect 1860 735 1890 740
rect 1860 715 1865 735
rect 1865 715 1885 735
rect 1885 715 1890 735
rect 1860 710 1890 715
rect 1860 635 1890 640
rect 1860 615 1865 635
rect 1865 615 1885 635
rect 1885 615 1890 635
rect 1860 610 1890 615
rect 1860 535 1890 540
rect 1860 515 1865 535
rect 1865 515 1885 535
rect 1885 515 1890 535
rect 1860 510 1890 515
rect 1860 435 1890 440
rect 1860 415 1865 435
rect 1865 415 1885 435
rect 1885 415 1890 435
rect 1860 410 1890 415
rect 1860 335 1890 340
rect 1860 315 1865 335
rect 1865 315 1885 335
rect 1885 315 1890 335
rect 1860 310 1890 315
rect 2060 635 2090 640
rect 2060 615 2065 635
rect 2065 615 2085 635
rect 2085 615 2090 635
rect 2060 610 2090 615
rect 2060 535 2090 540
rect 2060 515 2065 535
rect 2065 515 2085 535
rect 2085 515 2090 535
rect 2060 510 2090 515
rect 2060 435 2090 440
rect 2060 415 2065 435
rect 2065 415 2085 435
rect 2085 415 2090 435
rect 2060 410 2090 415
rect 2060 335 2090 340
rect 2060 315 2065 335
rect 2065 315 2085 335
rect 2085 315 2090 335
rect 2060 310 2090 315
rect 1860 210 1890 240
rect 1860 110 1890 140
rect 2460 635 2490 640
rect 2460 615 2465 635
rect 2465 615 2485 635
rect 2485 615 2490 635
rect 2460 610 2490 615
rect 2460 535 2490 540
rect 2460 515 2465 535
rect 2465 515 2485 535
rect 2485 515 2490 535
rect 2460 510 2490 515
rect 2460 435 2490 440
rect 2460 415 2465 435
rect 2465 415 2485 435
rect 2485 415 2490 435
rect 2460 410 2490 415
rect 2460 335 2490 340
rect 2460 315 2465 335
rect 2465 315 2485 335
rect 2485 315 2490 335
rect 2460 310 2490 315
rect 2060 210 2090 240
rect 2060 110 2090 140
rect 2660 735 2690 740
rect 2660 715 2665 735
rect 2665 715 2685 735
rect 2685 715 2690 735
rect 2660 710 2690 715
rect 2660 635 2690 640
rect 2660 615 2665 635
rect 2665 615 2685 635
rect 2685 615 2690 635
rect 2660 610 2690 615
rect 2660 535 2690 540
rect 2660 515 2665 535
rect 2665 515 2685 535
rect 2685 515 2690 535
rect 2660 510 2690 515
rect 2660 435 2690 440
rect 2660 415 2665 435
rect 2665 415 2685 435
rect 2685 415 2690 435
rect 2660 410 2690 415
rect 2660 335 2690 340
rect 2660 315 2665 335
rect 2665 315 2685 335
rect 2685 315 2690 335
rect 2660 310 2690 315
rect 2460 210 2490 240
rect 2460 110 2490 140
rect 2660 210 2690 240
rect 2660 110 2690 140
<< metal2 >>
rect 1450 3740 3100 3750
rect 1450 3710 1860 3740
rect 1890 3710 2060 3740
rect 2090 3710 2260 3740
rect 2290 3710 2460 3740
rect 2490 3710 2660 3740
rect 2690 3710 3100 3740
rect 1450 3700 3100 3710
rect 1450 3640 3100 3650
rect 1450 3610 1860 3640
rect 1890 3610 2060 3640
rect 2090 3610 2260 3640
rect 2290 3610 2460 3640
rect 2490 3610 2660 3640
rect 2690 3610 3100 3640
rect 1450 3600 3100 3610
rect 1450 3540 3100 3550
rect 1450 3510 1860 3540
rect 1890 3510 2060 3540
rect 2090 3510 2260 3540
rect 2290 3510 2460 3540
rect 2490 3510 2660 3540
rect 2690 3510 3100 3540
rect 1450 3500 3100 3510
rect 1450 3440 3100 3450
rect 1450 3410 1860 3440
rect 1890 3410 2060 3440
rect 2090 3410 2260 3440
rect 2290 3410 2460 3440
rect 2490 3410 2660 3440
rect 2690 3410 3100 3440
rect 1450 3400 3100 3410
rect 1450 3340 3100 3350
rect 1450 3310 1860 3340
rect 1890 3310 2060 3340
rect 2090 3310 2260 3340
rect 2290 3310 2460 3340
rect 2490 3310 2660 3340
rect 2690 3310 3100 3340
rect 1450 3300 3100 3310
rect 1450 3240 3100 3250
rect 1450 3210 1860 3240
rect 1890 3210 2060 3240
rect 2090 3210 2260 3240
rect 2290 3210 2460 3240
rect 2490 3210 2660 3240
rect 2690 3210 3100 3240
rect 1450 3200 3100 3210
rect 1450 3140 3100 3150
rect 1450 3110 1860 3140
rect 1890 3110 2060 3140
rect 2090 3110 2260 3140
rect 2290 3110 2460 3140
rect 2490 3110 2660 3140
rect 2690 3110 3100 3140
rect 1450 3100 3100 3110
rect 1950 3040 2000 3050
rect 1950 3010 1960 3040
rect 1990 3010 2000 3040
rect 1950 3000 2000 3010
rect 2150 3040 2200 3050
rect 2150 3010 2160 3040
rect 2190 3010 2200 3040
rect 2150 3000 2200 3010
rect 2350 3040 2400 3050
rect 2350 3010 2360 3040
rect 2390 3010 2400 3040
rect 2350 3000 2400 3010
rect 2550 3040 2600 3050
rect 2550 3010 2560 3040
rect 2590 3010 2600 3040
rect 2550 3000 2600 3010
rect 1450 2900 1850 2950
rect 2700 2900 3100 2950
rect 1450 2840 3100 2850
rect 1450 2810 1860 2840
rect 1890 2810 2060 2840
rect 2090 2810 2260 2840
rect 2290 2810 2460 2840
rect 2490 2810 2660 2840
rect 2690 2810 3100 2840
rect 1450 2800 3100 2810
rect 1450 2440 3100 2450
rect 1450 2410 1860 2440
rect 1890 2410 2260 2440
rect 2290 2410 2660 2440
rect 2690 2410 3100 2440
rect 1450 2400 3100 2410
rect 1450 2300 1850 2350
rect 2700 2300 3100 2350
rect 1450 2240 3100 2250
rect 1450 2210 1860 2240
rect 1890 2210 2260 2240
rect 2290 2210 2660 2240
rect 2690 2210 3100 2240
rect 1450 2200 3100 2210
rect 1450 2100 1850 2150
rect 2700 2100 3100 2150
rect 1450 2040 3100 2050
rect 1450 2010 1860 2040
rect 1890 2010 2260 2040
rect 2290 2010 2660 2040
rect 2690 2010 3100 2040
rect 1450 2000 3100 2010
rect 1950 1940 2000 1950
rect 1950 1910 1960 1940
rect 1990 1910 2000 1940
rect 1950 1900 2000 1910
rect 2150 1940 2200 1950
rect 2150 1910 2160 1940
rect 2190 1910 2200 1940
rect 2150 1900 2200 1910
rect 2350 1940 2400 1950
rect 2350 1910 2360 1940
rect 2390 1910 2400 1940
rect 2350 1900 2400 1910
rect 2550 1940 2600 1950
rect 2550 1910 2560 1940
rect 2590 1910 2600 1940
rect 2550 1900 2600 1910
rect 1450 1840 3100 1850
rect 1450 1810 1860 1840
rect 1890 1810 2260 1840
rect 2290 1810 2660 1840
rect 2690 1810 3100 1840
rect 1450 1800 3100 1810
rect 1450 1700 1850 1750
rect 2700 1700 3100 1750
rect 1450 1640 3100 1650
rect 1450 1610 1860 1640
rect 1890 1610 2260 1640
rect 2290 1610 2660 1640
rect 2690 1610 3100 1640
rect 1450 1600 3100 1610
rect 1450 1500 1850 1550
rect 2700 1500 3100 1550
rect 1450 1440 3100 1450
rect 1450 1410 1860 1440
rect 1890 1410 2260 1440
rect 2290 1410 2660 1440
rect 2690 1410 3100 1440
rect 1450 1400 3100 1410
rect 1450 1040 3100 1050
rect 1450 1010 1860 1040
rect 1890 1010 2060 1040
rect 2090 1010 2260 1040
rect 2290 1010 2460 1040
rect 2490 1010 2660 1040
rect 2690 1010 3100 1040
rect 1450 1000 3100 1010
rect 1450 900 1850 950
rect 2700 900 3100 950
rect 1950 840 2000 850
rect 1950 810 1960 840
rect 1990 810 2000 840
rect 1950 800 2000 810
rect 2150 840 2200 850
rect 2150 810 2160 840
rect 2190 810 2200 840
rect 2150 800 2200 810
rect 2350 840 2400 850
rect 2350 810 2360 840
rect 2390 810 2400 840
rect 2350 800 2400 810
rect 2550 840 2600 850
rect 2550 810 2560 840
rect 2590 810 2600 840
rect 2550 800 2600 810
rect 1450 740 3100 750
rect 1450 710 1860 740
rect 1890 710 2060 740
rect 2090 710 2260 740
rect 2290 710 2460 740
rect 2490 710 2660 740
rect 2690 710 3100 740
rect 1450 700 3100 710
rect 1450 640 3100 650
rect 1450 610 1860 640
rect 1890 610 2060 640
rect 2090 610 2260 640
rect 2290 610 2460 640
rect 2490 610 2660 640
rect 2690 610 3100 640
rect 1450 600 3100 610
rect 1950 550 2000 600
rect 2150 550 2200 600
rect 2350 550 2400 600
rect 2550 550 2600 600
rect 1450 540 3100 550
rect 1450 510 1860 540
rect 1890 510 2060 540
rect 2090 510 2260 540
rect 2290 510 2460 540
rect 2490 510 2660 540
rect 2690 510 3100 540
rect 1450 500 3100 510
rect 1950 450 2000 500
rect 2150 450 2200 500
rect 2350 450 2400 500
rect 2550 450 2600 500
rect 1450 440 3100 450
rect 1450 410 1860 440
rect 1890 410 2060 440
rect 2090 410 2260 440
rect 2290 410 2460 440
rect 2490 410 2660 440
rect 2690 410 3100 440
rect 1450 400 3100 410
rect 1950 350 2000 400
rect 2150 350 2200 400
rect 2350 350 2400 400
rect 2550 350 2600 400
rect 1450 340 3100 350
rect 1450 310 1860 340
rect 1890 310 2060 340
rect 2090 310 2260 340
rect 2290 310 2460 340
rect 2490 310 2660 340
rect 2690 310 3100 340
rect 1450 300 3100 310
rect 1950 250 2000 300
rect 2150 250 2200 300
rect 2350 250 2400 300
rect 2550 250 2600 300
rect 1450 240 3100 250
rect 1450 210 1860 240
rect 1890 210 2060 240
rect 2090 210 2260 240
rect 2290 210 2460 240
rect 2490 210 2660 240
rect 2690 210 3100 240
rect 1450 200 3100 210
rect 1450 140 3100 150
rect 1450 110 1860 140
rect 1890 110 2060 140
rect 2090 110 2260 140
rect 2290 110 2460 140
rect 2490 110 2660 140
rect 2690 110 3100 140
rect 1450 100 3100 110
<< via2 >>
rect 1860 3710 1890 3740
rect 2060 3710 2090 3740
rect 2260 3710 2290 3740
rect 2460 3710 2490 3740
rect 2660 3710 2690 3740
rect 1860 3610 1890 3640
rect 2060 3610 2090 3640
rect 2260 3610 2290 3640
rect 2460 3610 2490 3640
rect 2660 3610 2690 3640
rect 1860 3510 1890 3540
rect 2060 3510 2090 3540
rect 2260 3510 2290 3540
rect 2460 3510 2490 3540
rect 2660 3510 2690 3540
rect 1860 3410 1890 3440
rect 2060 3410 2090 3440
rect 2260 3410 2290 3440
rect 2460 3410 2490 3440
rect 2660 3410 2690 3440
rect 1860 3310 1890 3340
rect 2060 3310 2090 3340
rect 2260 3310 2290 3340
rect 2460 3310 2490 3340
rect 2660 3310 2690 3340
rect 1860 3210 1890 3240
rect 2060 3210 2090 3240
rect 2260 3210 2290 3240
rect 2460 3210 2490 3240
rect 2660 3210 2690 3240
rect 1860 3110 1890 3140
rect 2060 3110 2090 3140
rect 2260 3110 2290 3140
rect 2460 3110 2490 3140
rect 2660 3110 2690 3140
rect 1960 3010 1990 3040
rect 2160 3010 2190 3040
rect 2360 3010 2390 3040
rect 2560 3010 2590 3040
rect 1860 2810 1890 2840
rect 2060 2810 2090 2840
rect 2260 2810 2290 2840
rect 2460 2810 2490 2840
rect 2660 2810 2690 2840
rect 1860 2410 1890 2440
rect 2260 2410 2290 2440
rect 2660 2410 2690 2440
rect 1860 2210 1890 2240
rect 2260 2210 2290 2240
rect 2660 2210 2690 2240
rect 1860 2010 1890 2040
rect 2260 2010 2290 2040
rect 2660 2010 2690 2040
rect 1960 1910 1990 1940
rect 2160 1910 2190 1940
rect 2360 1910 2390 1940
rect 2560 1910 2590 1940
rect 1860 1810 1890 1840
rect 2260 1810 2290 1840
rect 2660 1810 2690 1840
rect 1860 1610 1890 1640
rect 2260 1610 2290 1640
rect 2660 1610 2690 1640
rect 1860 1410 1890 1440
rect 2260 1410 2290 1440
rect 2660 1410 2690 1440
rect 1860 1010 1890 1040
rect 2060 1010 2090 1040
rect 2260 1010 2290 1040
rect 2460 1010 2490 1040
rect 2660 1010 2690 1040
rect 1960 810 1990 840
rect 2160 810 2190 840
rect 2360 810 2390 840
rect 2560 810 2590 840
rect 1860 710 1890 740
rect 2060 710 2090 740
rect 2260 710 2290 740
rect 2460 710 2490 740
rect 2660 710 2690 740
rect 1860 610 1890 640
rect 2060 610 2090 640
rect 2260 610 2290 640
rect 2460 610 2490 640
rect 2660 610 2690 640
rect 1860 510 1890 540
rect 2060 510 2090 540
rect 2260 510 2290 540
rect 2460 510 2490 540
rect 2660 510 2690 540
rect 1860 410 1890 440
rect 2060 410 2090 440
rect 2260 410 2290 440
rect 2460 410 2490 440
rect 2660 410 2690 440
rect 1860 310 1890 340
rect 2060 310 2090 340
rect 2260 310 2290 340
rect 2460 310 2490 340
rect 2660 310 2690 340
rect 1860 210 1890 240
rect 2060 210 2090 240
rect 2260 210 2290 240
rect 2460 210 2490 240
rect 2660 210 2690 240
rect 1860 110 1890 140
rect 2060 110 2090 140
rect 2260 110 2290 140
rect 2460 110 2490 140
rect 2660 110 2690 140
<< metal3 >>
rect 1450 3740 3100 3750
rect 1450 3710 1860 3740
rect 1890 3710 2060 3740
rect 2090 3710 2260 3740
rect 2290 3710 2460 3740
rect 2490 3710 2660 3740
rect 2690 3710 3100 3740
rect 1450 3700 3100 3710
rect 1450 3640 3100 3650
rect 1450 3610 1860 3640
rect 1890 3610 2060 3640
rect 2090 3610 2260 3640
rect 2290 3610 2460 3640
rect 2490 3610 2660 3640
rect 2690 3610 3100 3640
rect 1450 3600 3100 3610
rect 1450 3540 3100 3550
rect 1450 3510 1860 3540
rect 1890 3510 2060 3540
rect 2090 3510 2260 3540
rect 2290 3510 2460 3540
rect 2490 3510 2660 3540
rect 2690 3510 3100 3540
rect 1450 3500 3100 3510
rect 1450 3440 3100 3450
rect 1450 3410 1860 3440
rect 1890 3410 2060 3440
rect 2090 3410 2260 3440
rect 2290 3410 2460 3440
rect 2490 3410 2660 3440
rect 2690 3410 3100 3440
rect 1450 3400 3100 3410
rect 1450 3340 3100 3350
rect 1450 3310 1860 3340
rect 1890 3310 2060 3340
rect 2090 3310 2260 3340
rect 2290 3310 2460 3340
rect 2490 3310 2660 3340
rect 2690 3310 3100 3340
rect 1450 3300 3100 3310
rect 1450 3240 3100 3250
rect 1450 3210 1860 3240
rect 1890 3210 2060 3240
rect 2090 3210 2260 3240
rect 2290 3210 2460 3240
rect 2490 3210 2660 3240
rect 2690 3210 3100 3240
rect 1450 3200 3100 3210
rect 1450 3140 3100 3150
rect 1450 3110 1860 3140
rect 1890 3110 2060 3140
rect 2090 3110 2260 3140
rect 2290 3110 2460 3140
rect 2490 3110 2660 3140
rect 2690 3110 3100 3140
rect 1450 3100 3100 3110
rect 1950 3045 2000 3050
rect 1950 3005 1955 3045
rect 1995 3005 2000 3045
rect 1950 3000 2000 3005
rect 2150 3045 2200 3050
rect 2150 3005 2155 3045
rect 2195 3005 2200 3045
rect 2150 3000 2200 3005
rect 2350 3045 2400 3050
rect 2350 3005 2355 3045
rect 2395 3005 2400 3045
rect 2350 3000 2400 3005
rect 2550 3045 2600 3050
rect 2550 3005 2555 3045
rect 2595 3005 2600 3045
rect 2550 3000 2600 3005
rect 1450 2900 1850 2950
rect 2700 2900 3100 2950
rect 1450 2840 3100 2850
rect 1450 2810 1860 2840
rect 1890 2810 2060 2840
rect 2090 2810 2260 2840
rect 2290 2810 2460 2840
rect 2490 2810 2660 2840
rect 2690 2810 3100 2840
rect 1450 2800 3100 2810
rect 1450 2440 3100 2450
rect 1450 2410 1860 2440
rect 1890 2410 2260 2440
rect 2290 2410 2660 2440
rect 2690 2410 3100 2440
rect 1450 2400 3100 2410
rect 1450 2240 3100 2250
rect 1450 2210 1860 2240
rect 1890 2210 2260 2240
rect 2290 2210 2660 2240
rect 2690 2210 3100 2240
rect 1450 2200 3100 2210
rect 1450 2040 3100 2050
rect 1450 2010 1860 2040
rect 1890 2010 2260 2040
rect 2290 2010 2660 2040
rect 2690 2010 3100 2040
rect 1450 2000 3100 2010
rect 1950 1945 2000 1950
rect 1950 1905 1955 1945
rect 1995 1905 2000 1945
rect 1950 1900 2000 1905
rect 2150 1945 2200 1950
rect 2150 1905 2155 1945
rect 2195 1905 2200 1945
rect 2150 1900 2200 1905
rect 2350 1945 2400 1950
rect 2350 1905 2355 1945
rect 2395 1905 2400 1945
rect 2350 1900 2400 1905
rect 2550 1945 2600 1950
rect 2550 1905 2555 1945
rect 2595 1905 2600 1945
rect 2550 1900 2600 1905
rect 1450 1840 3100 1850
rect 1450 1810 1860 1840
rect 1890 1810 2260 1840
rect 2290 1810 2660 1840
rect 2690 1810 3100 1840
rect 1450 1800 3100 1810
rect 1450 1745 3100 1750
rect 1450 1705 1955 1745
rect 1995 1705 2555 1745
rect 2595 1705 3100 1745
rect 1450 1700 3100 1705
rect 1450 1640 3100 1650
rect 1450 1610 1860 1640
rect 1890 1610 2260 1640
rect 2290 1610 2660 1640
rect 2690 1610 3100 1640
rect 1450 1600 3100 1610
rect 1450 1440 3100 1450
rect 1450 1410 1860 1440
rect 1890 1410 2260 1440
rect 2290 1410 2660 1440
rect 2690 1410 3100 1440
rect 1450 1400 3100 1410
rect 1450 1040 3100 1050
rect 1450 1010 1860 1040
rect 1890 1010 2060 1040
rect 2090 1010 2260 1040
rect 2290 1010 2460 1040
rect 2490 1010 2660 1040
rect 2690 1010 3100 1040
rect 1450 1000 3100 1010
rect 1450 900 1850 950
rect 2700 900 3100 950
rect 1950 845 2000 850
rect 1950 805 1955 845
rect 1995 805 2000 845
rect 1950 800 2000 805
rect 2150 845 2200 850
rect 2150 805 2155 845
rect 2195 805 2200 845
rect 2150 800 2200 805
rect 2350 845 2400 850
rect 2350 805 2355 845
rect 2395 805 2400 845
rect 2350 800 2400 805
rect 2550 845 2600 850
rect 2550 805 2555 845
rect 2595 805 2600 845
rect 2550 800 2600 805
rect 1450 740 3100 750
rect 1450 710 1860 740
rect 1890 710 2060 740
rect 2090 710 2260 740
rect 2290 710 2460 740
rect 2490 710 2660 740
rect 2690 710 3100 740
rect 1450 700 3100 710
rect 1450 640 3100 650
rect 1450 610 1860 640
rect 1890 610 2060 640
rect 2090 610 2260 640
rect 2290 610 2460 640
rect 2490 610 2660 640
rect 2690 610 3100 640
rect 1450 600 3100 610
rect 1950 550 2000 600
rect 2150 550 2200 600
rect 2350 550 2400 600
rect 2550 550 2600 600
rect 1450 540 3100 550
rect 1450 510 1860 540
rect 1890 510 2060 540
rect 2090 510 2260 540
rect 2290 510 2460 540
rect 2490 510 2660 540
rect 2690 510 3100 540
rect 1450 500 3100 510
rect 1950 450 2000 500
rect 2150 450 2200 500
rect 2350 450 2400 500
rect 2550 450 2600 500
rect 1450 440 3100 450
rect 1450 410 1860 440
rect 1890 410 2060 440
rect 2090 410 2260 440
rect 2290 410 2460 440
rect 2490 410 2660 440
rect 2690 410 3100 440
rect 1450 400 3100 410
rect 1950 350 2000 400
rect 2150 350 2200 400
rect 2350 350 2400 400
rect 2550 350 2600 400
rect 1450 340 3100 350
rect 1450 310 1860 340
rect 1890 310 2060 340
rect 2090 310 2260 340
rect 2290 310 2460 340
rect 2490 310 2660 340
rect 2690 310 3100 340
rect 1450 300 3100 310
rect 1950 250 2000 300
rect 2150 250 2200 300
rect 2350 250 2400 300
rect 2550 250 2600 300
rect 1450 240 3100 250
rect 1450 210 1860 240
rect 1890 210 2060 240
rect 2090 210 2260 240
rect 2290 210 2460 240
rect 2490 210 2660 240
rect 2690 210 3100 240
rect 1450 200 3100 210
rect 1450 140 3100 150
rect 1450 110 1860 140
rect 1890 110 2060 140
rect 2090 110 2260 140
rect 2290 110 2460 140
rect 2490 110 2660 140
rect 2690 110 3100 140
rect 1450 100 3100 110
<< via3 >>
rect 1955 3040 1995 3045
rect 1955 3010 1960 3040
rect 1960 3010 1990 3040
rect 1990 3010 1995 3040
rect 1955 3005 1995 3010
rect 2155 3040 2195 3045
rect 2155 3010 2160 3040
rect 2160 3010 2190 3040
rect 2190 3010 2195 3040
rect 2155 3005 2195 3010
rect 2355 3040 2395 3045
rect 2355 3010 2360 3040
rect 2360 3010 2390 3040
rect 2390 3010 2395 3040
rect 2355 3005 2395 3010
rect 2555 3040 2595 3045
rect 2555 3010 2560 3040
rect 2560 3010 2590 3040
rect 2590 3010 2595 3040
rect 2555 3005 2595 3010
rect 1955 1940 1995 1945
rect 1955 1910 1960 1940
rect 1960 1910 1990 1940
rect 1990 1910 1995 1940
rect 1955 1905 1995 1910
rect 2155 1940 2195 1945
rect 2155 1910 2160 1940
rect 2160 1910 2190 1940
rect 2190 1910 2195 1940
rect 2155 1905 2195 1910
rect 2355 1940 2395 1945
rect 2355 1910 2360 1940
rect 2360 1910 2390 1940
rect 2390 1910 2395 1940
rect 2355 1905 2395 1910
rect 2555 1940 2595 1945
rect 2555 1910 2560 1940
rect 2560 1910 2590 1940
rect 2590 1910 2595 1940
rect 2555 1905 2595 1910
rect 1955 1705 1995 1745
rect 2555 1705 2595 1745
rect 1955 840 1995 845
rect 1955 810 1960 840
rect 1960 810 1990 840
rect 1990 810 1995 840
rect 1955 805 1995 810
rect 2155 840 2195 845
rect 2155 810 2160 840
rect 2160 810 2190 840
rect 2190 810 2195 840
rect 2155 805 2195 810
rect 2355 840 2395 845
rect 2355 810 2360 840
rect 2360 810 2390 840
rect 2390 810 2395 840
rect 2355 805 2395 810
rect 2555 840 2595 845
rect 2555 810 2560 840
rect 2560 810 2590 840
rect 2590 810 2595 840
rect 2555 805 2595 810
<< metal4 >>
rect 1950 3045 2000 3050
rect 1950 3005 1955 3045
rect 1995 3005 2000 3045
rect 1950 1945 2000 3005
rect 1950 1905 1955 1945
rect 1995 1905 2000 1945
rect 1950 1745 2000 1905
rect 1950 1705 1955 1745
rect 1995 1705 2000 1745
rect 1950 845 2000 1705
rect 1950 805 1955 845
rect 1995 805 2000 845
rect 1950 800 2000 805
rect 2150 3045 2200 3050
rect 2150 3005 2155 3045
rect 2195 3005 2200 3045
rect 2150 1945 2200 3005
rect 2150 1905 2155 1945
rect 2195 1905 2200 1945
rect 2150 845 2200 1905
rect 2150 805 2155 845
rect 2195 805 2200 845
rect 2150 800 2200 805
rect 2350 3045 2400 3050
rect 2350 3005 2355 3045
rect 2395 3005 2400 3045
rect 2350 1945 2400 3005
rect 2350 1905 2355 1945
rect 2395 1905 2400 1945
rect 2350 845 2400 1905
rect 2350 805 2355 845
rect 2395 805 2400 845
rect 2350 800 2400 805
rect 2550 3045 2600 3050
rect 2550 3005 2555 3045
rect 2595 3005 2600 3045
rect 2550 1945 2600 3005
rect 2550 1905 2555 1945
rect 2595 1905 2600 1945
rect 2550 1745 2600 1905
rect 2550 1705 2555 1745
rect 2595 1705 2600 1745
rect 2550 845 2600 1705
rect 2550 805 2555 845
rect 2595 805 2600 845
rect 2550 800 2600 805
<< labels >>
rlabel metal3 1450 1700 3100 1750 0 ref
port 1 nsew
rlabel metal1 2050 1900 2100 1950 0 x
rlabel locali 1750 3650 2800 3700 0 bp
port 2 nsew
rlabel locali 1750 2750 2800 2800 0 bn
port 3 nsew
rlabel metal3 1450 3700 3100 3750 0 vdd
port 4 nsew
rlabel metal3 1450 100 3100 150 0 vdd
port 4 nsew
rlabel metal3 1450 2800 3100 2850 0 vss
port 5 nsew
rlabel metal3 1450 1000 3100 1050 0 vss
port 5 nsew
<< end >>
